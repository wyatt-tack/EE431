magic
tech sky130A
timestamp 1729544331
<< nwell >>
rect 1130 700 1350 960
<< nmos >>
rect 1210 610 1250 660
<< pmos >>
rect 1210 720 1250 820
<< ndiff >>
rect 1170 650 1210 660
rect 1170 620 1180 650
rect 1200 620 1210 650
rect 1170 610 1210 620
rect 1250 650 1290 660
rect 1250 620 1260 650
rect 1280 620 1290 650
rect 1250 610 1290 620
<< pdiff >>
rect 1150 810 1210 820
rect 1150 730 1160 810
rect 1200 730 1210 810
rect 1150 720 1210 730
rect 1250 810 1310 820
rect 1250 730 1260 810
rect 1300 730 1310 810
rect 1250 720 1310 730
<< ndiffc >>
rect 1180 620 1200 650
rect 1260 620 1280 650
<< pdiffc >>
rect 1160 730 1200 810
rect 1260 730 1300 810
<< psubdiff >>
rect 1150 550 1310 570
rect 1150 530 1170 550
rect 1290 530 1310 550
rect 1150 510 1310 530
<< nsubdiff >>
rect 1150 910 1330 930
rect 1150 880 1170 910
rect 1310 880 1330 910
rect 1150 860 1330 880
<< psubdiffcont >>
rect 1170 530 1290 550
<< nsubdiffcont >>
rect 1170 880 1310 910
<< poly >>
rect 1210 820 1250 840
rect 1210 660 1250 720
rect 1210 590 1250 610
<< locali >>
rect 1150 910 1330 930
rect 1150 880 1170 910
rect 1310 880 1330 910
rect 1150 860 1330 880
rect 1150 820 1190 860
rect 1150 810 1210 820
rect 1150 730 1160 810
rect 1200 730 1210 810
rect 1150 720 1210 730
rect 1250 810 1310 820
rect 1250 730 1260 810
rect 1300 730 1310 810
rect 1250 720 1310 730
rect 1250 660 1280 720
rect 1170 650 1210 660
rect 1170 620 1180 650
rect 1200 620 1210 650
rect 1170 610 1210 620
rect 1250 650 1290 660
rect 1250 620 1260 650
rect 1280 620 1290 650
rect 1250 610 1290 620
rect 1170 570 1200 610
rect 1150 550 1310 570
rect 1150 530 1170 550
rect 1290 530 1310 550
rect 1150 510 1310 530
<< viali >>
rect 1170 880 1310 910
rect 1170 530 1290 550
<< metal1 >>
rect 1080 910 1400 940
rect 1080 880 1170 910
rect 1310 880 1400 910
rect 1080 850 1400 880
rect 1080 550 1400 580
rect 1080 530 1170 550
rect 1290 530 1400 550
rect 1080 500 1400 530
<< end >>
