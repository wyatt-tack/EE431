* NGSPICE file created from pwm.ext - technology: sky130A

.subckt magic_nand A B Y VDD VSS a_100_n230#
X0 Y A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.5 pd=2.5 as=0.9 ps=4.9 w=2 l=0.5
**devattr s=36000,980 d=20000,500
X1 Y B a_100_n230# VSS sky130_fd_pr__nfet_01v8 ad=0.9 pd=4.9 as=0.5 ps=2.5 w=2 l=0.5
**devattr s=20000,500 d=36000,980
X2 a_100_n230# A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.5 pd=2.5 as=0.9 ps=4.9 w=2 l=0.5
**devattr s=36000,980 d=20000,500
X3 VDD B Y VDD sky130_fd_pr__pfet_01v8 ad=0.9 pd=4.9 as=0.5 ps=2.5 w=2 l=0.5
**devattr s=20000,500 d=36000,980
C0 Y A 0.09013f
C1 B a_100_n230# 0.014208f
C2 B Y 0.253425f
C3 Y a_100_n230# 0.017664f
C4 VDD A 0.202433f
C5 B VDD 0.118732f
C6 a_100_n230# VDD 0.002196f
C7 Y VDD 0.207993f
C8 B A 0.21018f
C9 Y VSS 0.271727f
C10 B VSS 0.476474f
C11 A VSS 0.453547f
C12 VDD VSS 1.23585f
C13 a_100_n230# VSS 0.028228f
.ends

.subckt magic_inv X Y VDD VSS
X0 Y X VDD VDD sky130_fd_pr__pfet_01v8 ad=0.9 pd=4.9 as=0.9 ps=4.9 w=2 l=0.5
**devattr s=36000,980 d=36000,980
X1 Y X VSS VSS sky130_fd_pr__nfet_01v8 ad=0.45 pd=2.9 as=0.45 ps=2.9 w=1 l=0.5
**devattr s=18000,580 d=18000,580
C0 VDD X 0.197978f
C1 Y X 0.105971f
C2 VDD Y 0.10691f
C3 Y VSS 0.267668f
C4 X VSS 0.481952f
C5 VDD VSS 0.843976f
.ends

.subckt magic_dff clk Q magic_nand_2/Y magic_nand_3/Y notQ magic_nand_1/a_100_n230#
+ magic_nand_2/a_100_n230# magic_inv_0/Y D VDD VSS
Xmagic_nand_0 magic_nand_3/Y notQ Q VDD VSS magic_nand_0/a_100_n230# magic_nand
Xmagic_nand_1 Q magic_nand_2/Y notQ VDD VSS magic_nand_1/a_100_n230# magic_nand
Xmagic_nand_2 magic_inv_0/Y clk magic_nand_2/Y VDD VSS magic_nand_2/a_100_n230# magic_nand
Xmagic_nand_3 clk D magic_nand_3/Y VDD VSS magic_nand_3/a_100_n230# magic_nand
Xmagic_inv_0 D magic_inv_0/Y VDD VSS magic_inv
C0 magic_nand_3/Y clk 5.03e-19
C1 Q magic_nand_2/Y 0.070054f
C2 magic_nand_3/Y D 0.013145f
C3 magic_nand_2/Y magic_nand_3/a_100_n230# 0.003027f
C4 magic_nand_3/Y notQ 0.112791f
C5 VDD magic_nand_2/Y 0.013097f
C6 Q clk 0.022129f
C7 Q D 3.91e-19
C8 Q magic_inv_0/Y 3.16e-19
C9 magic_nand_3/a_100_n230# clk 9.29e-20
C10 Q notQ 0.204136f
C11 magic_nand_3/a_100_n230# D 6.62e-20
C12 VDD clk 0.276198f
C13 VDD D 0.282719f
C14 VDD magic_inv_0/Y 0.082291f
C15 Q magic_nand_3/Y 0.011129f
C16 VDD notQ 0.444233f
C17 VDD magic_nand_0/a_100_n230# 0.009399f
C18 magic_nand_2/Y clk 0.005838f
C19 magic_nand_2/Y D 0.005584f
C20 magic_nand_2/Y magic_inv_0/Y 0.005014f
C21 VDD magic_nand_3/Y 0.06714f
C22 magic_nand_2/Y notQ 0.027101f
C23 magic_nand_2/a_100_n230# clk 3.18e-19
C24 magic_nand_2/Y magic_nand_1/a_100_n230# 1.53e-19
C25 clk D 0.512204f
C26 magic_nand_2/Y magic_nand_3/Y 0.003303f
C27 magic_inv_0/Y clk 0.126572f
C28 magic_inv_0/Y D 0.025042f
C29 clk notQ 6.78e-19
C30 VDD Q 0.780984f
C31 notQ D 0.004634f
C32 VDD magic_nand_3/a_100_n230# 0.007823f
C33 magic_nand_0/a_100_n230# notQ 0.008218f
C34 VDD VSS 6.870138f
C35 D VSS 1.396145f
C36 magic_nand_3/Y VSS 0.626503f
C37 magic_nand_3/a_100_n230# VSS 0.028228f
C38 magic_nand_2/Y VSS 0.830572f
C39 clk VSS 3.249527f
C40 magic_inv_0/Y VSS 0.560832f
C41 magic_nand_2/a_100_n230# VSS 0.040303f
C42 Q VSS 1.533211f
C43 magic_nand_1/a_100_n230# VSS 0.034833f
C44 notQ VSS 1.445663f
C45 magic_nand_0/a_100_n230# VSS 0.028228f
.ends

.subckt magic_xnor A magic_nand_1/Y magic_nand_2/Y magic_nand_1/a_100_n230# magic_nand_0/a_100_n230#
+ magic_inv_1/Y magic_nand_2/a_100_n230# magic_inv_0/Y B VDD Y VSS
Xmagic_nand_0 magic_nand_1/Y magic_nand_2/Y Y VDD VSS magic_nand_0/a_100_n230# magic_nand
Xmagic_nand_1 A B magic_nand_1/Y VDD VSS magic_nand_1/a_100_n230# magic_nand
Xmagic_nand_2 magic_inv_0/Y magic_inv_1/Y magic_nand_2/Y VDD VSS magic_nand_2/a_100_n230#
+ magic_nand
Xmagic_inv_0 B magic_inv_0/Y VDD VSS magic_inv
Xmagic_inv_1 A magic_inv_1/Y VDD VSS magic_inv
C0 Y VDD 0.016266f
C1 VSS magic_nand_2/a_100_n230# 0.012357f
C2 magic_nand_0/a_100_n230# magic_inv_1/Y 1.14e-19
C3 magic_inv_0/Y magic_inv_1/Y 0.134093f
C4 Y B 3.91e-19
C5 Y magic_nand_2/Y 0.074699f
C6 B VDD 0.134682f
C7 VDD magic_nand_2/Y 0.072046f
C8 B magic_nand_2/Y 0.002564f
C9 VSS Y -0.029084f
C10 VSS VDD 0.742841f
C11 VSS B 0.023906f
C12 VSS magic_nand_2/Y 0.190942f
C13 Y magic_nand_0/a_100_n230# -0.013335f
C14 magic_nand_0/a_100_n230# VDD -0.001132f
C15 magic_nand_1/Y magic_inv_1/Y 2.81e-19
C16 magic_inv_0/Y VDD 0.082312f
C17 magic_nand_0/a_100_n230# magic_nand_2/Y 0.038774f
C18 B magic_inv_0/Y 0.015802f
C19 magic_inv_0/Y magic_nand_2/Y 0.016464f
C20 magic_nand_1/a_100_n230# magic_inv_1/Y 1.71e-19
C21 VSS magic_nand_0/a_100_n230# -0.022613f
C22 VSS magic_inv_0/Y 0.027978f
C23 A magic_inv_1/Y 0.01498f
C24 Y magic_nand_1/Y -0.005512f
C25 magic_nand_1/Y VDD 0.02847f
C26 magic_inv_1/Y magic_nand_2/a_100_n230# 3.18e-19
C27 B magic_nand_1/Y 0.015962f
C28 magic_nand_1/Y magic_nand_2/Y 0.07956f
C29 magic_nand_1/a_100_n230# VDD 0.009875f
C30 Y magic_inv_1/Y 2.91e-19
C31 VSS magic_nand_1/Y 0.083428f
C32 magic_inv_1/Y VDD 0.073805f
C33 A VDD 0.242512f
C34 magic_nand_1/a_100_n230# B 1.42e-19
C35 B magic_inv_1/Y 0.051559f
C36 magic_inv_1/Y magic_nand_2/Y 0.021402f
C37 A B 0.175283f
C38 A magic_nand_2/Y 6e-19
C39 magic_nand_0/a_100_n230# magic_nand_1/Y 3.07e-20
C40 magic_nand_1/Y magic_inv_0/Y 0.021701f
C41 VSS magic_inv_1/Y 0.464243f
C42 VSS A 0.04505f
C43 VDD 0 5.241346f
C44 VSS 0 -0.106448f
C45 magic_nand_2/Y 0 0.735869f
C46 magic_inv_1/Y 0 0.876545f
C47 magic_inv_0/Y 0 0.513873f
C48 magic_nand_2/a_100_n230# 0 0.028228f
C49 magic_nand_1/Y 0 0.570102f
C50 B 0 0.998797f
C51 A 0 1.186725f
C52 magic_nand_1/a_100_n230# 0 0.028228f
C53 Y 0 0.299583f
C54 magic_nand_0/a_100_n230# 0 0.028228f
.ends

.subckt magic_and A Y VDD B magic_nand_0/a_100_n230# magic_inv_0/X VSS
Xmagic_nand_0 A B magic_inv_0/X VDD VSS magic_nand_0/a_100_n230# magic_nand
Xmagic_inv_0 magic_inv_0/X Y VDD VSS magic_inv
C0 VDD magic_inv_0/X 0.005293f
C1 VDD Y 0.001742f
C2 magic_inv_0/X VSS 0.09428f
C3 VSS A 0.003964f
C4 magic_nand_0/a_100_n230# VSS 0.004912f
C5 magic_inv_0/X B 0.013119f
C6 Y B 4.88e-19
C7 VDD B 0.005182f
C8 B VSS 0.009819f
C9 Y magic_inv_0/X 0.010551f
C10 VSS 0 3.79e-20
C11 Y 0 0.252201f
C12 VDD 0 1.901415f
C13 magic_inv_0/X 0 0.650359f
C14 B 0 0.460323f
C15 A 0 0.453547f
C16 magic_nand_0/a_100_n230# 0 0.028228f
.ends

.subckt magic_comp A0 A1 Y magic_and_1/magic_inv_0/X magic_and_1/B magic_xnor_1/magic_inv_1/Y
+ magic_xnor_1/magic_inv_0/Y magic_xnor_0/magic_nand_2/Y magic_xnor_2/magic_nand_1/Y
+ magic_and_2/magic_inv_0/X magic_xnor_2/magic_inv_0/Y magic_xnor_2/magic_inv_1/Y
+ magic_xnor_3/magic_nand_1/Y A3 magic_xnor_1/magic_nand_2/Y magic_and_0/B magic_xnor_3/magic_nand_0/a_100_n230#
+ B0 magic_xnor_3/magic_nand_2/Y magic_xnor_3/magic_nand_1/a_100_n230# magic_and_2/B
+ magic_xnor_3/magic_inv_1/Y B3 magic_and_1/A magic_xnor_0/magic_nand_1/Y magic_xnor_3/magic_inv_0/Y
+ magic_xnor_2/magic_nand_2/Y magic_and_0/magic_inv_0/X magic_and_0/A magic_xnor_0/magic_inv_1/Y
+ magic_xnor_0/magic_inv_0/Y VDD B1 A2 magic_and_2/A magic_xnor_1/magic_nand_1/Y VSS
+ B2
Xmagic_xnor_0 B0 magic_xnor_0/magic_nand_1/Y magic_xnor_0/magic_nand_2/Y magic_xnor_0/magic_nand_1/a_100_n230#
+ magic_xnor_0/magic_nand_0/a_100_n230# magic_xnor_0/magic_inv_1/Y magic_xnor_0/magic_nand_2/a_100_n230#
+ magic_xnor_0/magic_inv_0/Y A0 VDD magic_and_0/B VSS magic_xnor
Xmagic_xnor_1 B1 magic_xnor_1/magic_nand_1/Y magic_xnor_1/magic_nand_2/Y magic_xnor_1/magic_nand_1/a_100_n230#
+ magic_xnor_1/magic_nand_0/a_100_n230# magic_xnor_1/magic_inv_1/Y magic_xnor_1/magic_nand_2/a_100_n230#
+ magic_xnor_1/magic_inv_0/Y A1 VDD magic_and_0/A VSS magic_xnor
Xmagic_xnor_2 B2 magic_xnor_2/magic_nand_1/Y magic_xnor_2/magic_nand_2/Y magic_xnor_2/magic_nand_1/a_100_n230#
+ magic_xnor_2/magic_nand_0/a_100_n230# magic_xnor_2/magic_inv_1/Y magic_xnor_2/magic_nand_2/a_100_n230#
+ magic_xnor_2/magic_inv_0/Y A2 VDD magic_and_1/A VSS magic_xnor
Xmagic_xnor_3 B3 magic_xnor_3/magic_nand_1/Y magic_xnor_3/magic_nand_2/Y magic_xnor_3/magic_nand_1/a_100_n230#
+ magic_xnor_3/magic_nand_0/a_100_n230# magic_xnor_3/magic_inv_1/Y magic_xnor_3/magic_nand_2/a_100_n230#
+ magic_xnor_3/magic_inv_0/Y A3 VDD magic_and_2/A VSS magic_xnor
Xmagic_and_0 magic_and_0/A magic_and_1/B VDD magic_and_0/B magic_and_0/magic_nand_0/a_100_n230#
+ magic_and_0/magic_inv_0/X VSS magic_and
Xmagic_and_1 magic_and_1/A magic_and_2/B VDD magic_and_1/B magic_and_1/magic_nand_0/a_100_n230#
+ magic_and_1/magic_inv_0/X VSS magic_and
Xmagic_and_2 magic_and_2/A Y VDD magic_and_2/B magic_and_2/magic_nand_0/a_100_n230#
+ magic_and_2/magic_inv_0/X VSS magic_and
C0 A3 A2 1.739336f
C1 magic_and_0/B VSS 0.322655f
C2 magic_and_0/B magic_xnor_0/magic_inv_1/Y 0.004862f
C3 magic_xnor_2/magic_inv_1/Y magic_and_1/B 0.001122f
C4 B1 magic_xnor_1/magic_nand_1/Y 6.29e-19
C5 magic_and_1/magic_inv_0/X magic_xnor_2/magic_inv_0/Y 7.57e-19
C6 VSS magic_and_1/magic_inv_0/X 0.00493f
C7 magic_xnor_1/magic_inv_1/Y magic_and_1/B 7.65e-20
C8 magic_and_2/magic_inv_0/X A3 0.001223f
C9 B0 VDD 0.217725f
C10 magic_xnor_1/magic_nand_1/Y A1 0.002948f
C11 magic_and_1/magic_inv_0/X magic_and_2/A 0.003363f
C12 B2 VDD 0.458517f
C13 VSS magic_xnor_0/magic_inv_0/Y 3.91e-20
C14 magic_and_0/magic_inv_0/X magic_xnor_1/magic_nand_1/Y 3.43e-20
C15 magic_and_0/magic_inv_0/X magic_and_1/A 0.003363f
C16 magic_and_0/B magic_xnor_1/magic_inv_1/Y 0.01381f
C17 magic_xnor_2/magic_inv_1/Y magic_and_1/magic_inv_0/X 6.54e-19
C18 magic_and_1/magic_inv_0/X magic_xnor_2/magic_nand_1/Y 3.43e-20
C19 magic_and_1/magic_nand_0/a_100_n230# magic_and_1/B 3.05e-20
C20 magic_and_0/A magic_xnor_2/magic_nand_2/Y 9.88e-19
C21 magic_and_0/A magic_xnor_1/magic_nand_2/Y 0.157912f
C22 magic_and_0/A A2 0.085823f
C23 B2 A3 0.032768f
C24 magic_and_0/magic_inv_0/X magic_xnor_1/magic_inv_0/Y 7.57e-19
C25 magic_and_2/B magic_and_1/magic_inv_0/X 0.00375f
C26 VDD magic_xnor_3/magic_nand_1/Y 0.001607f
C27 VDD magic_xnor_3/magic_nand_2/Y 6.99e-19
C28 VSS magic_xnor_3/magic_inv_1/Y 0.065528f
C29 magic_and_2/A magic_xnor_3/magic_inv_1/Y 0.116308f
C30 VDD magic_xnor_2/magic_inv_0/Y 8.48e-19
C31 VDD VSS 2.22109f
C32 VDD magic_xnor_0/magic_inv_1/Y 0.015491f
C33 VDD magic_and_2/A 0.512407f
C34 magic_and_0/B B1 0.020686f
C35 magic_xnor_2/magic_inv_1/Y magic_xnor_3/magic_inv_1/Y 3.28e-20
C36 magic_xnor_1/magic_nand_2/Y A2 0.011525f
C37 magic_and_0/magic_inv_0/X magic_and_1/B 0.00375f
C38 VDD magic_xnor_0/magic_nand_2/a_100_n230# 3.88e-19
C39 magic_and_0/B A1 0.093186f
C40 Y magic_and_2/magic_inv_0/X 0.002706f
C41 B0 magic_xnor_0/magic_nand_2/Y 1.93e-19
C42 magic_xnor_2/magic_inv_1/Y VDD 0.001633f
C43 VDD magic_xnor_2/magic_nand_1/Y 0.005274f
C44 magic_and_0/magic_inv_0/X magic_and_0/B 0.001364f
C45 B0 A0 0.041536f
C46 B1 magic_xnor_0/magic_inv_0/Y 5.27e-20
C47 A3 magic_xnor_3/magic_nand_1/Y 0.002948f
C48 VDD magic_xnor_1/magic_inv_1/Y 0.001633f
C49 VDD B3 0.332265f
C50 B2 A0 0.034392f
C51 B2 magic_and_0/A 0.016031f
C52 magic_and_1/A magic_xnor_3/magic_inv_0/Y 9.2e-20
C53 magic_and_0/magic_inv_0/X magic_and_1/magic_inv_0/X 7.26e-21
C54 A3 VSS 0.003625f
C55 magic_and_2/B magic_xnor_3/magic_inv_1/Y 0.001122f
C56 A3 magic_and_2/A 4.36e-19
C57 magic_and_2/B VDD 0.004945f
C58 VDD magic_xnor_1/magic_nand_0/a_100_n230# 6.22e-19
C59 magic_and_1/A magic_and_1/B 0.061618f
C60 A3 magic_xnor_2/magic_nand_1/Y 0.022873f
C61 VDD magic_xnor_2/magic_nand_0/a_100_n230# 6.22e-19
C62 B2 magic_xnor_1/magic_nand_2/Y 0.020436f
C63 B2 A2 0.486209f
C64 A3 B3 0.700245f
C65 magic_and_0/B magic_xnor_1/magic_nand_1/a_100_n230# 5.94e-20
C66 magic_and_0/B magic_xnor_1/magic_nand_1/Y 0.001166f
C67 magic_xnor_0/magic_nand_2/Y VSS -0.006408f
C68 B1 VDD 0.617586f
C69 magic_and_1/A magic_and_1/magic_inv_0/X 0.046398f
C70 magic_and_0/A magic_xnor_2/magic_inv_0/Y 9.2e-20
C71 VSS A0 7.9e-19
C72 magic_xnor_3/magic_nand_2/a_100_n230# VSS 1.59e-19
C73 magic_and_0/A VSS 0.560822f
C74 VDD A1 0.78035f
C75 magic_xnor_3/magic_nand_2/a_100_n230# magic_and_2/A 0.008718f
C76 magic_xnor_0/magic_nand_1/Y VDD 0.004772f
C77 magic_xnor_1/magic_nand_2/a_100_n230# magic_and_0/A 0.008718f
C78 magic_xnor_1/magic_inv_0/Y magic_and_1/B 9.81e-20
C79 magic_and_0/magic_inv_0/X VDD 0.002386f
C80 magic_xnor_2/magic_inv_1/Y magic_and_0/A 0.012688f
C81 magic_xnor_1/magic_inv_0/Y magic_and_0/B 9.2e-20
C82 magic_and_0/A magic_xnor_2/magic_nand_1/Y 0.001166f
C83 A0 B3 0.080192f
C84 magic_and_0/A magic_xnor_1/magic_inv_1/Y 0.116308f
C85 B0 B2 0.018364f
C86 Y VSS 0.116668f
C87 magic_xnor_1/magic_nand_2/Y magic_xnor_2/magic_inv_0/Y 3.03e-21
C88 VSS magic_xnor_2/magic_nand_2/Y -0.006235f
C89 Y magic_and_2/A 0.048107f
C90 magic_xnor_1/magic_nand_2/Y VSS -0.006235f
C91 VSS A2 0.003673f
C92 magic_and_2/magic_inv_0/X magic_xnor_3/magic_nand_1/Y 3.43e-20
C93 magic_and_0/B magic_and_1/B 2.03e-24
C94 magic_and_2/magic_inv_0/X VSS 0.034941f
C95 magic_and_1/A magic_xnor_3/magic_inv_1/Y 0.012688f
C96 magic_and_2/magic_inv_0/X magic_and_2/A 0.046398f
C97 magic_xnor_1/magic_nand_1/a_100_n230# VDD 6.99e-19
C98 magic_and_1/magic_inv_0/X magic_and_1/B 0.001566f
C99 A2 magic_xnor_2/magic_nand_1/Y 0.002948f
C100 B3 magic_xnor_2/magic_nand_2/Y 0.015825f
C101 VDD magic_xnor_1/magic_nand_1/Y 0.004688f
C102 magic_and_1/A VDD 0.637375f
C103 A2 B3 0.102095f
C104 magic_xnor_0/magic_nand_2/Y B1 0.041193f
C105 magic_and_2/magic_inv_0/X B3 2.93e-19
C106 magic_and_0/B magic_xnor_0/magic_inv_0/Y 2.6e-19
C107 VDD magic_xnor_2/magic_nand_1/a_100_n230# 6.99e-19
C108 B1 A0 0.064621f
C109 magic_xnor_0/magic_nand_2/Y A1 0.017422f
C110 magic_and_0/A B1 0.009691f
C111 A0 A1 0.107301f
C112 B0 VSS 0.031873f
C113 magic_and_0/A A1 4.36e-19
C114 B2 VSS 0.019736f
C115 magic_xnor_1/magic_inv_0/Y VDD 8.48e-19
C116 magic_and_0/magic_inv_0/X magic_and_0/A 0.046398f
C117 magic_and_1/A A3 0.081673f
C118 magic_and_2/magic_inv_0/X magic_and_2/B 0.001566f
C119 B2 magic_xnor_2/magic_nand_1/Y 6.29e-19
C120 B0 B3 6.28e-19
C121 B2 magic_xnor_1/magic_inv_1/Y 0.005651f
C122 B1 A2 0.036498f
C123 B2 B3 1.6929f
C124 VDD magic_and_1/B 0.004945f
C125 A2 A1 1.014962f
C126 magic_and_0/B VDD 0.207216f
C127 VSS magic_xnor_3/magic_nand_2/Y -0.006249f
C128 magic_and_2/A magic_xnor_3/magic_nand_2/Y 0.157912f
C129 VDD magic_and_1/magic_inv_0/X 0.002386f
C130 VSS magic_xnor_2/magic_inv_0/Y 0.002448f
C131 magic_and_1/A magic_and_0/A 0.006892f
C132 magic_and_2/magic_nand_0/a_100_n230# VSS 0.001392f
C133 magic_xnor_0/magic_inv_1/Y VSS 0.062078f
C134 VDD magic_xnor_0/magic_inv_0/Y 0.004118f
C135 VSS magic_and_2/A 0.543962f
C136 magic_xnor_1/magic_nand_2/a_100_n230# VSS 1.59e-19
C137 B3 magic_xnor_3/magic_nand_1/Y 6.29e-19
C138 VDD magic_xnor_0/magic_nand_1/a_100_n230# 6.99e-19
C139 magic_and_0/A magic_xnor_2/magic_nand_1/a_100_n230# 5.94e-20
C140 magic_xnor_2/magic_inv_1/Y VSS 0.065676f
C141 B0 B1 0.415585f
C142 B2 B1 1.076414f
C143 magic_xnor_1/magic_inv_1/Y magic_xnor_2/magic_inv_0/Y 1.15e-20
C144 magic_xnor_1/magic_inv_0/Y magic_xnor_0/magic_nand_2/Y 3.03e-21
C145 B3 magic_xnor_2/magic_inv_0/Y 1.67e-20
C146 VSS magic_xnor_1/magic_inv_1/Y 0.065676f
C147 B0 A1 0.050185f
C148 VSS B3 0.018158f
C149 magic_xnor_0/magic_inv_1/Y magic_xnor_1/magic_inv_1/Y 3.28e-20
C150 B2 A1 0.132649f
C151 magic_xnor_0/magic_nand_1/Y B0 8.29e-19
C152 magic_and_1/A magic_xnor_2/magic_nand_2/Y 0.157912f
C153 magic_and_2/A B3 0.009691f
C154 magic_xnor_1/magic_nand_1/Y A2 0.029803f
C155 magic_xnor_0/magic_nand_1/Y B2 2.61e-19
C156 magic_and_1/A A2 4.36e-19
C157 magic_xnor_1/magic_inv_0/Y magic_and_0/A 0.012015f
C158 magic_xnor_2/magic_inv_1/Y magic_xnor_1/magic_inv_1/Y 3.28e-20
C159 magic_xnor_2/magic_inv_1/Y B3 0.005651f
C160 magic_xnor_2/magic_nand_1/Y B3 0.011024f
C161 magic_and_2/B magic_xnor_2/magic_inv_0/Y 9.81e-20
C162 magic_and_2/magic_nand_0/a_100_n230# magic_and_2/B 3.05e-20
C163 magic_and_2/B VSS 0.01737f
C164 VSS magic_and_1/magic_nand_0/a_100_n230# 2.17e-19
C165 magic_and_2/B magic_and_2/A 0.061619f
C166 VSS magic_xnor_2/magic_nand_2/a_100_n230# 1.59e-19
C167 magic_and_0/A magic_and_1/B 0.043537f
C168 Y magic_xnor_3/magic_inv_0/Y 1.24e-19
C169 magic_xnor_0/magic_nand_0/a_100_n230# VDD 6.22e-19
C170 magic_xnor_3/magic_inv_0/Y magic_xnor_2/magic_nand_2/Y 3.03e-21
C171 magic_and_0/B magic_xnor_0/magic_nand_2/Y 0.141165f
C172 magic_xnor_2/magic_inv_1/Y magic_and_2/B 7.65e-20
C173 magic_and_0/B A0 1.17e-19
C174 magic_and_0/B magic_and_0/A 0.158653f
C175 magic_and_2/B B3 0.001222f
C176 magic_and_2/magic_inv_0/X magic_xnor_3/magic_inv_0/Y 7.57e-19
C177 B1 VSS 0.023016f
C178 B1 magic_xnor_0/magic_inv_1/Y 0.005651f
C179 B2 magic_xnor_1/magic_nand_1/Y 0.017161f
C180 A3 magic_xnor_3/magic_inv_1/Y 1.42e-32
C181 B2 magic_and_1/A 0.009691f
C182 VSS A1 0.003673f
C183 magic_and_0/magic_inv_0/X VSS 0.004879f
C184 VDD A3 1.162519f
C185 magic_and_0/B magic_xnor_1/magic_nand_2/Y 9.88e-19
C186 B1 B3 0.001349f
C187 B3 A1 0.09995f
C188 magic_and_1/magic_inv_0/X A2 0.001223f
C189 magic_xnor_0/magic_nand_1/Y B3 9.75e-20
C190 magic_and_0/magic_inv_0/X magic_xnor_1/magic_inv_1/Y 6.54e-19
C191 B2 magic_xnor_1/magic_inv_0/Y 3.57e-20
C192 magic_and_2/magic_inv_0/X magic_and_1/magic_inv_0/X 7.26e-21
C193 magic_and_1/A magic_xnor_3/magic_nand_1/Y 0.001166f
C194 magic_and_1/A magic_xnor_3/magic_nand_2/Y 9.88e-19
C195 magic_xnor_0/magic_nand_2/Y VDD 0.008234f
C196 magic_and_1/A magic_xnor_3/magic_nand_1/a_100_n230# 5.94e-20
C197 magic_and_1/A magic_xnor_2/magic_inv_0/Y 0.012015f
C198 VDD A0 0.061379f
C199 magic_and_0/A VDD 0.629023f
C200 magic_and_1/A VSS 0.561339f
C201 B2 magic_and_1/B 0.001222f
C202 magic_and_1/A magic_and_2/A 0.006892f
C203 B0 magic_and_0/B 2.5e-19
C204 magic_and_1/A magic_xnor_2/magic_inv_1/Y 0.116308f
C205 Y magic_xnor_3/magic_inv_1/Y 9.91e-20
C206 B1 A1 0.306032f
C207 B2 magic_and_1/magic_inv_0/X 2.93e-19
C208 magic_xnor_0/magic_nand_1/Y B1 0.042386f
C209 magic_and_1/A B3 0.014558f
C210 magic_and_0/magic_inv_0/X B1 2.93e-19
C211 VDD magic_xnor_2/magic_nand_2/Y 0.007048f
C212 magic_xnor_3/magic_inv_0/Y VSS 0.003026f
C213 magic_xnor_0/magic_nand_1/Y A1 0.044988f
C214 magic_xnor_1/magic_nand_2/Y VDD 0.006794f
C215 VDD A2 0.944114f
C216 magic_xnor_1/magic_inv_0/Y VSS 0.002448f
C217 magic_xnor_3/magic_inv_0/Y magic_and_2/A 0.012015f
C218 magic_xnor_1/magic_inv_0/Y magic_xnor_0/magic_inv_1/Y 1.15e-20
C219 magic_and_0/magic_inv_0/X A1 0.001223f
C220 magic_and_2/magic_inv_0/X magic_xnor_3/magic_inv_1/Y 6.54e-19
C221 magic_and_2/magic_inv_0/X VDD 8.33e-19
C222 magic_xnor_2/magic_inv_1/Y magic_xnor_3/magic_inv_0/Y 1.15e-20
C223 magic_and_1/A magic_and_2/B 0.043537f
C224 magic_and_1/A magic_xnor_2/magic_nand_2/a_100_n230# 0.008718f
C225 VSS magic_and_1/B 0.011683f
C226 A3 magic_xnor_2/magic_nand_2/Y 0.00868f
C227 Y 0 0.539191f
C228 magic_and_2/magic_inv_0/X 0 0.650359f
C229 magic_and_2/B 0 1.005271f
C230 magic_and_2/magic_nand_0/a_100_n230# 0 0.028228f
C231 magic_and_1/magic_inv_0/X 0 0.650359f
C232 magic_and_1/B 0 1.005271f
C233 magic_and_1/magic_nand_0/a_100_n230# 0 0.028228f
C234 VDD 0 26.95971f
C235 magic_and_0/magic_inv_0/X 0 0.650359f
C236 magic_and_0/magic_nand_0/a_100_n230# 0 0.028228f
C237 magic_xnor_3/magic_nand_2/Y 0 0.735869f
C238 magic_xnor_3/magic_inv_1/Y 0 0.876545f
C239 magic_xnor_3/magic_inv_0/Y 0 0.513873f
C240 magic_xnor_3/magic_nand_2/a_100_n230# 0 0.028228f
C241 magic_xnor_3/magic_nand_1/Y 0 0.570102f
C242 A3 0 1.833927f
C243 B3 0 3.097305f
C244 magic_xnor_3/magic_nand_1/a_100_n230# 0 0.028228f
C245 magic_and_2/A 0 1.742389f
C246 magic_xnor_3/magic_nand_0/a_100_n230# 0 0.028228f
C247 magic_xnor_2/magic_nand_2/Y 0 0.735869f
C248 magic_xnor_2/magic_inv_1/Y 0 0.876545f
C249 magic_xnor_2/magic_inv_0/Y 0 0.513873f
C250 magic_xnor_2/magic_nand_2/a_100_n230# 0 0.028228f
C251 magic_xnor_2/magic_nand_1/Y 0 0.570102f
C252 A2 0 1.444479f
C253 B2 0 2.326525f
C254 magic_xnor_2/magic_nand_1/a_100_n230# 0 0.028228f
C255 magic_and_1/A 0 1.548071f
C256 magic_xnor_2/magic_nand_0/a_100_n230# 0 0.028228f
C257 VSS 0 0.155042f
C258 magic_xnor_1/magic_nand_2/Y 0 0.735869f
C259 magic_xnor_1/magic_inv_1/Y 0 0.876545f
C260 magic_xnor_1/magic_inv_0/Y 0 0.513873f
C261 magic_xnor_1/magic_nand_2/a_100_n230# 0 0.028228f
C262 magic_xnor_1/magic_nand_1/Y 0 0.570102f
C263 A1 0 1.401717f
C264 B1 0 2.835861f
C265 magic_xnor_1/magic_nand_1/a_100_n230# 0 0.028228f
C266 magic_and_0/A 0 1.481641f
C267 magic_xnor_1/magic_nand_0/a_100_n230# 0 0.028228f
C268 magic_xnor_0/magic_nand_2/Y 0 0.735869f
C269 magic_xnor_0/magic_inv_1/Y 0 0.876545f
C270 magic_xnor_0/magic_inv_0/Y 0 0.513873f
C271 magic_xnor_0/magic_nand_2/a_100_n230# 0 0.028228f
C272 magic_xnor_0/magic_nand_1/Y 0 0.570102f
C273 A0 0 0.982813f
C274 B0 0 1.769344f
C275 magic_xnor_0/magic_nand_1/a_100_n230# 0 0.028228f
C276 magic_and_0/B 0 1.359748f
C277 magic_xnor_0/magic_nand_0/a_100_n230# 0 0.028228f
.ends

.subckt magic_etdff clk magic_dff_1/magic_nand_1/a_100_n230# magic_dff_0/magic_nand_3/Y
+ magic_dff_1/magic_nand_2/a_100_n230# magic_dff_0/magic_inv_0/Y magic_dff_1/magic_nand_3/Y
+ notQ magic_inv_1/Y magic_dff_1/magic_inv_0/Y magic_dff_0/magic_nand_2/Y magic_dff_1/D
+ magic_inv_1/X magic_dff_0/notQ D magic_dff_1/magic_nand_2/Y VDD Q VSS
Xmagic_dff_0 magic_inv_1/X magic_dff_1/D magic_dff_0/magic_nand_2/Y magic_dff_0/magic_nand_3/Y
+ magic_dff_0/notQ magic_dff_0/magic_nand_1/a_100_n230# magic_dff_0/magic_nand_2/a_100_n230#
+ magic_dff_0/magic_inv_0/Y D VDD VSS magic_dff
Xmagic_dff_1 magic_inv_1/Y Q magic_dff_1/magic_nand_2/Y magic_dff_1/magic_nand_3/Y
+ notQ magic_dff_1/magic_nand_1/a_100_n230# magic_dff_1/magic_nand_2/a_100_n230# magic_dff_1/magic_inv_0/Y
+ magic_dff_1/D VDD VSS magic_dff
Xmagic_inv_0 clk magic_inv_1/X VDD VSS magic_inv
Xmagic_inv_1 magic_inv_1/X magic_inv_1/Y VDD VSS magic_inv
C0 magic_inv_1/Y magic_dff_0/magic_nand_1/a_100_n230# 0.008718f
C1 magic_dff_0/magic_nand_3/Y magic_dff_1/D 1.26e-19
C2 magic_inv_1/Y magic_dff_0/magic_inv_0/Y 0.017008f
C3 magic_dff_0/notQ magic_inv_1/Y 0.083427f
C4 clk VDD 0.009114f
C5 magic_inv_1/Y VDD 0.062853f
C6 magic_inv_1/X clk 0.021739f
C7 magic_inv_1/Y magic_inv_1/X 0.260754f
C8 magic_inv_1/Y magic_dff_1/magic_inv_0/Y 2.6e-20
C9 magic_dff_0/magic_nand_2/Y magic_inv_1/Y 0.061361f
C10 magic_dff_0/notQ VDD 7.2e-19
C11 magic_dff_1/D magic_inv_1/Y 0.082207f
C12 magic_dff_0/notQ magic_dff_1/magic_inv_0/Y 0.003242f
C13 notQ VDD 1.06e-19
C14 magic_dff_0/notQ magic_dff_1/magic_nand_3/Y 6.01e-20
C15 VDD Q 0.00382f
C16 notQ Q 9.94e-19
C17 magic_dff_1/magic_nand_2/Y notQ 2.15e-19
C18 magic_inv_1/X VDD 0.339081f
C19 magic_dff_1/magic_nand_3/Y VDD 2.12e-19
C20 D clk 0.023212f
C21 D magic_inv_1/Y 0.084411f
C22 magic_dff_0/notQ magic_dff_1/D 0.08104f
C23 magic_dff_0/magic_nand_2/Y magic_dff_1/magic_inv_0/Y 4.14e-19
C24 magic_dff_1/D VDD 0.050093f
C25 magic_dff_0/magic_nand_3/Y magic_inv_1/Y 1.59e-19
C26 magic_dff_1/D magic_dff_1/magic_nand_3/Y 0.001872f
C27 magic_dff_0/magic_nand_2/Y magic_dff_1/D 1.04e-20
C28 D VDD 0.123858f
C29 D magic_inv_1/X 0.100784f
C30 magic_dff_0/magic_nand_3/Y VDD 7.84e-20
C31 magic_inv_1/Y magic_dff_0/magic_nand_2/a_100_n230# 0.008718f
C32 magic_dff_0/magic_nand_3/Y magic_inv_1/X 0.002282f
C33 magic_inv_1/X VSS 3.219988f
C34 clk VSS 0.513302f
C35 VDD VSS 14.160234f
C36 magic_dff_1/D VSS 2.570121f
C37 magic_dff_1/magic_nand_3/Y VSS 0.625399f
C38 magic_dff_1/magic_nand_3/a_100_n230# VSS 0.028228f
C39 magic_dff_1/magic_nand_2/Y VSS 0.670071f
C40 magic_inv_1/Y VSS 4.860871f
C41 magic_dff_1/magic_inv_0/Y VSS 0.538833f
C42 magic_dff_1/magic_nand_2/a_100_n230# VSS 0.028228f
C43 Q VSS 1.439376f
C44 magic_dff_1/magic_nand_1/a_100_n230# VSS 0.028228f
C45 notQ VSS 1.098129f
C46 magic_dff_1/magic_nand_0/a_100_n230# VSS 0.028228f
C47 D VSS 1.527642f
C48 magic_dff_0/magic_nand_3/Y VSS 0.625399f
C49 magic_dff_0/magic_nand_3/a_100_n230# VSS 0.028228f
C50 magic_dff_0/magic_nand_2/Y VSS 0.66738f
C51 magic_dff_0/magic_inv_0/Y VSS 0.539688f
C52 magic_dff_0/magic_nand_2/a_100_n230# VSS 0.028578f
C53 magic_dff_0/magic_nand_1/a_100_n230# VSS 0.029266f
C54 magic_dff_0/notQ VSS 1.079399f
C55 magic_dff_0/magic_nand_0/a_100_n230# VSS 0.028228f
.ends

.subckt magic_counter clk S0 S1 S2 S3 magic_etdff_1/magic_dff_1/D magic_etdff_0/magic_dff_1/magic_nand_3/Y
+ magic_etdff_3/magic_dff_1/magic_nand_2/Y magic_etdff_2/magic_dff_0/notQ magic_etdff_1/magic_inv_1/Y
+ magic_etdff_1/magic_dff_1/magic_nand_3/Y magic_etdff_2/magic_dff_0/magic_inv_0/Y
+ magic_etdff_3/magic_dff_1/magic_nand_1/a_100_n230# magic_etdff_2/magic_dff_1/D magic_etdff_1/magic_inv_1/X
+ magic_etdff_3/magic_dff_0/magic_inv_0/Y magic_etdff_1/magic_dff_0/notQ magic_etdff_2/magic_dff_1/magic_inv_0/Y
+ magic_etdff_3/magic_dff_1/magic_nand_3/Y magic_etdff_2/magic_dff_0/magic_nand_2/Y
+ magic_etdff_0/D magic_etdff_0/magic_inv_1/Y magic_etdff_0/magic_dff_1/D magic_etdff_0/magic_inv_1/X
+ magic_etdff_3/magic_dff_0/notQ magic_etdff_2/D magic_etdff_3/magic_dff_1/magic_inv_0/Y
+ magic_etdff_0/magic_dff_0/magic_nand_3/Y magic_etdff_3/magic_inv_1/X magic_etdff_3/magic_inv_1/Y
+ magic_etdff_3/magic_dff_0/magic_nand_2/Y magic_etdff_2/magic_inv_1/X magic_etdff_1/D
+ magic_etdff_0/magic_dff_0/notQ magic_etdff_2/magic_dff_1/magic_nand_2/Y magic_etdff_0/magic_dff_0/magic_inv_0/Y
+ magic_etdff_3/magic_dff_1/D magic_etdff_1/magic_dff_0/magic_nand_3/Y VSS magic_etdff_3/D
+ VDD magic_etdff_2/magic_inv_1/Y
Xmagic_etdff_0 clk magic_etdff_0/magic_dff_1/magic_nand_1/a_100_n230# magic_etdff_0/magic_dff_0/magic_nand_3/Y
+ magic_etdff_0/magic_dff_1/magic_nand_2/a_100_n230# magic_etdff_0/magic_dff_0/magic_inv_0/Y
+ magic_etdff_0/magic_dff_1/magic_nand_3/Y magic_etdff_0/D magic_etdff_0/magic_inv_1/Y
+ magic_etdff_0/magic_dff_1/magic_inv_0/Y magic_etdff_0/magic_dff_0/magic_nand_2/Y
+ magic_etdff_0/magic_dff_1/D magic_etdff_0/magic_inv_1/X magic_etdff_0/magic_dff_0/notQ
+ magic_etdff_0/D magic_etdff_0/magic_dff_1/magic_nand_2/Y VDD S0 VSS magic_etdff
Xmagic_etdff_1 S0 magic_etdff_1/magic_dff_1/magic_nand_1/a_100_n230# magic_etdff_1/magic_dff_0/magic_nand_3/Y
+ magic_etdff_1/magic_dff_1/magic_nand_2/a_100_n230# magic_etdff_1/magic_dff_0/magic_inv_0/Y
+ magic_etdff_1/magic_dff_1/magic_nand_3/Y magic_etdff_1/D magic_etdff_1/magic_inv_1/Y
+ magic_etdff_1/magic_dff_1/magic_inv_0/Y magic_etdff_1/magic_dff_0/magic_nand_2/Y
+ magic_etdff_1/magic_dff_1/D magic_etdff_1/magic_inv_1/X magic_etdff_1/magic_dff_0/notQ
+ magic_etdff_1/D magic_etdff_1/magic_dff_1/magic_nand_2/Y VDD S1 VSS magic_etdff
Xmagic_etdff_2 S1 magic_etdff_2/magic_dff_1/magic_nand_1/a_100_n230# magic_etdff_2/magic_dff_0/magic_nand_3/Y
+ magic_etdff_2/magic_dff_1/magic_nand_2/a_100_n230# magic_etdff_2/magic_dff_0/magic_inv_0/Y
+ magic_etdff_2/magic_dff_1/magic_nand_3/Y magic_etdff_2/D magic_etdff_2/magic_inv_1/Y
+ magic_etdff_2/magic_dff_1/magic_inv_0/Y magic_etdff_2/magic_dff_0/magic_nand_2/Y
+ magic_etdff_2/magic_dff_1/D magic_etdff_2/magic_inv_1/X magic_etdff_2/magic_dff_0/notQ
+ magic_etdff_2/D magic_etdff_2/magic_dff_1/magic_nand_2/Y VDD S2 VSS magic_etdff
Xmagic_etdff_3 S2 magic_etdff_3/magic_dff_1/magic_nand_1/a_100_n230# magic_etdff_3/magic_dff_0/magic_nand_3/Y
+ magic_etdff_3/magic_dff_1/magic_nand_2/a_100_n230# magic_etdff_3/magic_dff_0/magic_inv_0/Y
+ magic_etdff_3/magic_dff_1/magic_nand_3/Y magic_etdff_3/D magic_etdff_3/magic_inv_1/Y
+ magic_etdff_3/magic_dff_1/magic_inv_0/Y magic_etdff_3/magic_dff_0/magic_nand_2/Y
+ magic_etdff_3/magic_dff_1/D magic_etdff_3/magic_inv_1/X magic_etdff_3/magic_dff_0/notQ
+ magic_etdff_3/D magic_etdff_3/magic_dff_1/magic_nand_2/Y VDD S3 VSS magic_etdff
C0 magic_etdff_3/magic_inv_1/X VDD 0.006701f
C1 magic_etdff_0/magic_dff_1/magic_inv_0/Y S1 4.78e-19
C2 magic_etdff_2/magic_dff_0/notQ magic_etdff_0/D 8.03e-19
C3 magic_etdff_2/magic_dff_0/magic_nand_3/Y magic_etdff_0/magic_dff_1/D 0.004383f
C4 magic_etdff_2/D magic_etdff_0/D 0.001606f
C5 magic_etdff_0/D magic_etdff_0/magic_dff_1/D 0.001408f
C6 S2 magic_etdff_0/D 1.25e-19
C7 magic_etdff_0/magic_dff_1/magic_inv_0/Y VDD 0.001022f
C8 magic_etdff_2/D magic_etdff_3/D 0.125665f
C9 S2 magic_etdff_3/D 0.075506f
C10 magic_etdff_1/magic_dff_1/magic_nand_1/a_100_n230# magic_etdff_1/D 0.00545f
C11 magic_etdff_2/magic_dff_0/magic_nand_3/Y magic_etdff_0/magic_inv_1/Y 4.9e-19
C12 S1 VDD 1.363633f
C13 S1 magic_etdff_3/magic_dff_1/magic_nand_3/Y 0.014898f
C14 magic_etdff_3/magic_dff_0/magic_nand_2/Y S2 4.7e-20
C15 magic_etdff_0/D magic_etdff_0/magic_inv_1/Y 1.006191f
C16 VDD magic_etdff_2/magic_dff_1/magic_nand_2/Y 4.92e-19
C17 magic_etdff_1/magic_dff_0/magic_inv_0/Y S0 0.01029f
C18 S0 magic_etdff_2/D 6.32e-21
C19 S0 S2 1.20837f
C20 magic_etdff_3/magic_inv_1/Y S2 0.058461f
C21 S1 magic_etdff_2/magic_inv_1/X 0.030211f
C22 magic_etdff_0/D magic_etdff_2/magic_inv_1/Y 0.001608f
C23 magic_etdff_2/magic_inv_1/X VDD 1.57e-19
C24 magic_etdff_0/D magic_etdff_0/magic_dff_0/magic_inv_0/Y 8.75e-19
C25 S1 magic_etdff_0/magic_inv_1/X 0.003922f
C26 S3 S2 0.020942f
C27 magic_etdff_1/magic_dff_0/magic_inv_0/Y magic_etdff_1/D 3.3e-19
C28 magic_etdff_2/magic_dff_1/D magic_etdff_2/D 0.001336f
C29 S0 magic_etdff_1/magic_dff_0/magic_nand_2/Y 0.009909f
C30 clk VDD 0.002002f
C31 magic_etdff_0/magic_inv_1/X VDD 0.001553f
C32 magic_etdff_0/magic_dff_1/magic_nand_2/Y magic_etdff_0/D 0.036891f
C33 magic_etdff_0/magic_dff_0/magic_nand_2/Y magic_etdff_2/magic_dff_0/magic_nand_3/Y 2.01e-20
C34 magic_etdff_3/magic_dff_0/notQ S2 0.032829f
C35 magic_etdff_2/magic_inv_1/X magic_etdff_0/magic_inv_1/X 0.001257f
C36 magic_etdff_2/magic_dff_1/D magic_etdff_0/magic_inv_1/Y 0.003587f
C37 magic_etdff_0/magic_dff_0/magic_nand_2/Y magic_etdff_0/D 8.03e-19
C38 magic_etdff_2/magic_dff_1/magic_nand_3/Y magic_etdff_0/D 8.85e-19
C39 magic_etdff_3/magic_dff_1/magic_nand_2/Y magic_etdff_3/D 0.035472f
C40 magic_etdff_1/magic_dff_0/magic_nand_2/Y magic_etdff_1/D 3.07e-19
C41 magic_etdff_2/magic_dff_1/magic_nand_1/a_100_n230# magic_etdff_2/D 0.005219f
C42 magic_etdff_2/magic_dff_1/magic_nand_3/Y magic_etdff_3/D 8.1e-20
C43 S0 magic_etdff_0/magic_dff_1/magic_nand_2/Y 0.008298f
C44 S0 magic_etdff_1/magic_dff_1/magic_nand_3/Y 1.75e-19
C45 magic_etdff_3/magic_inv_1/X magic_etdff_2/D 0.001672f
C46 magic_etdff_1/magic_dff_1/magic_nand_1/a_100_n230# VDD 0.004571f
C47 magic_etdff_3/magic_inv_1/X S2 0.08124f
C48 S0 magic_etdff_2/magic_dff_1/magic_nand_3/Y 0.004383f
C49 magic_etdff_2/magic_dff_0/notQ S1 0.002567f
C50 S1 magic_etdff_2/D 0.0064f
C51 magic_etdff_3/magic_dff_1/magic_inv_0/Y magic_etdff_3/D 0.005944f
C52 magic_etdff_3/D magic_etdff_3/magic_dff_1/D 0.001336f
C53 S1 magic_etdff_0/magic_dff_1/D 8.88e-19
C54 S2 S1 0.724876f
C55 magic_etdff_2/D magic_etdff_2/magic_dff_1/magic_nand_2/Y 0.035472f
C56 magic_etdff_1/magic_inv_1/X magic_etdff_0/D 9.29e-20
C57 S0 magic_etdff_1/magic_dff_0/magic_nand_3/Y 2.66e-21
C58 VDD magic_etdff_2/D 0.08532f
C59 VDD magic_etdff_0/magic_dff_1/D 0.002781f
C60 S2 VDD 1.12582f
C61 S2 magic_etdff_3/magic_dff_1/magic_nand_3/Y 0.043613f
C62 S0 magic_etdff_0/magic_dff_1/magic_nand_3/Y 1.14e-19
C63 S1 magic_etdff_0/magic_inv_1/Y 4.85e-19
C64 magic_etdff_2/magic_inv_1/X magic_etdff_2/D 0.027311f
C65 magic_etdff_2/D magic_etdff_2/magic_dff_0/magic_nand_2/Y 7.48e-19
C66 S0 magic_etdff_1/magic_inv_1/X 0.082068f
C67 magic_etdff_0/magic_dff_1/magic_inv_0/Y magic_etdff_2/magic_inv_1/Y 0.004524f
C68 VDD magic_etdff_0/magic_inv_1/Y 4.4e-19
C69 magic_etdff_0/magic_inv_1/X magic_etdff_2/D 0.003478f
C70 S1 magic_etdff_2/magic_inv_1/Y 0.018275f
C71 S1 magic_etdff_0/magic_dff_0/magic_inv_0/Y 4.78e-19
C72 S0 magic_etdff_1/magic_dff_1/magic_inv_0/Y 0.009868f
C73 magic_etdff_2/magic_inv_1/X magic_etdff_0/magic_inv_1/Y 0.001067f
C74 magic_etdff_0/magic_dff_1/magic_nand_3/Y magic_etdff_1/D 7.72e-20
C75 S0 magic_etdff_1/magic_dff_1/magic_nand_2/Y 0.020897f
C76 magic_etdff_3/D magic_etdff_3/magic_dff_0/magic_inv_0/Y 8.18e-19
C77 magic_etdff_0/magic_dff_1/magic_nand_1/a_100_n230# magic_etdff_0/D 0.00545f
C78 VDD magic_etdff_2/magic_inv_1/Y 1.5e-19
C79 VDD magic_etdff_0/magic_dff_0/magic_inv_0/Y 0.001022f
C80 magic_etdff_2/magic_dff_0/magic_nand_3/Y magic_etdff_0/D 8.85e-19
C81 magic_etdff_1/magic_inv_1/X magic_etdff_1/D 0.027773f
C82 S1 magic_etdff_0/magic_dff_1/magic_nand_2/Y 4.27e-19
C83 S0 magic_etdff_1/magic_inv_1/Y 0.086733f
C84 S1 magic_etdff_1/magic_dff_1/magic_nand_3/Y 1.43e-19
C85 magic_etdff_2/magic_inv_1/X magic_etdff_0/magic_dff_0/magic_inv_0/Y 0.004524f
C86 magic_etdff_1/magic_dff_1/magic_inv_0/Y magic_etdff_1/D 0.005753f
C87 magic_etdff_0/magic_dff_0/magic_nand_2/Y S1 4.27e-19
C88 magic_etdff_1/magic_dff_1/magic_nand_2/Y magic_etdff_1/D 0.036395f
C89 magic_etdff_2/magic_dff_1/magic_nand_3/Y S1 0.016845f
C90 magic_etdff_0/magic_dff_1/magic_nand_2/Y VDD 3.84e-19
C91 S0 magic_etdff_0/D 0.025107f
C92 magic_etdff_3/magic_dff_0/magic_nand_3/Y S1 0.014898f
C93 magic_etdff_3/magic_dff_0/magic_nand_2/Y magic_etdff_3/D 7.48e-19
C94 magic_etdff_0/magic_dff_0/magic_nand_2/Y VDD 3.84e-19
C95 magic_etdff_1/D magic_etdff_1/magic_inv_1/Y 1.00689f
C96 magic_etdff_3/magic_inv_1/Y magic_etdff_3/D 0.88731f
C97 magic_etdff_0/D magic_etdff_0/magic_dff_1/magic_nand_2/a_100_n230# 0.00545f
C98 magic_etdff_2/magic_dff_1/D magic_etdff_0/D 9.28e-19
C99 magic_etdff_1/D magic_etdff_0/D 0.116931f
C100 S1 magic_etdff_3/magic_dff_1/D 0.014319f
C101 S3 magic_etdff_3/D 0.007057f
C102 magic_etdff_2/magic_dff_0/notQ magic_etdff_0/magic_dff_1/D 6.32e-21
C103 S2 magic_etdff_2/D 0.012523f
C104 magic_etdff_2/magic_dff_1/magic_inv_0/Y magic_etdff_2/D 0.005944f
C105 S0 S3 3.6e-19
C106 magic_etdff_2/magic_dff_0/notQ magic_etdff_0/magic_inv_1/Y 4.27e-19
C107 S0 magic_etdff_1/D 1.02558f
C108 magic_etdff_2/D magic_etdff_0/magic_inv_1/Y 4.27e-19
C109 magic_etdff_2/D magic_etdff_2/magic_dff_0/magic_inv_0/Y 8.18e-19
C110 magic_etdff_1/magic_inv_1/X VDD 0.003295f
C111 magic_etdff_1/magic_dff_1/magic_nand_2/Y S1 9.55e-19
C112 magic_etdff_1/magic_dff_1/magic_nand_2/Y VDD 0.016199f
C113 magic_etdff_2/D magic_etdff_2/magic_dff_1/magic_nand_2/a_100_n230# 0.005219f
C114 magic_etdff_2/D magic_etdff_2/magic_inv_1/Y 0.88731f
C115 magic_etdff_1/D magic_etdff_1/magic_dff_1/magic_nand_2/a_100_n230# 0.00545f
C116 magic_etdff_0/magic_dff_1/D magic_etdff_2/magic_inv_1/Y 0.001585f
C117 magic_etdff_3/magic_inv_1/X magic_etdff_3/D 0.027311f
C118 magic_etdff_0/magic_dff_1/magic_inv_0/Y magic_etdff_0/D 0.006291f
C119 magic_etdff_2/magic_dff_0/magic_nand_3/Y S1 0.016845f
C120 magic_etdff_0/magic_inv_1/Y magic_etdff_2/magic_inv_1/Y 0.001407f
C121 magic_etdff_0/magic_dff_1/magic_nand_2/Y magic_etdff_2/D 0.003478f
C122 S1 magic_etdff_0/D 1.913593f
C123 magic_etdff_3/magic_dff_1/magic_nand_2/a_100_n230# magic_etdff_3/D 0.005219f
C124 magic_etdff_2/magic_dff_0/notQ magic_etdff_0/magic_dff_0/magic_nand_2/Y 0.003478f
C125 S1 magic_etdff_3/D 0.003187f
C126 magic_etdff_3/magic_dff_1/magic_nand_2/Y S2 4.7e-20
C127 magic_etdff_3/D magic_etdff_2/magic_dff_1/magic_nand_2/Y 4.26e-19
C128 VDD magic_etdff_0/D 0.194434f
C129 magic_etdff_2/magic_dff_1/magic_nand_3/Y S2 1.13e-19
C130 VDD magic_etdff_3/D 0.089509f
C131 S0 magic_etdff_1/magic_dff_0/notQ 0.002477f
C132 S0 S1 0.711168f
C133 magic_etdff_3/magic_inv_1/Y S1 0.015351f
C134 magic_etdff_3/magic_dff_0/magic_nand_3/Y S2 0.043724f
C135 magic_etdff_2/magic_inv_1/X magic_etdff_0/D 0.003931f
C136 magic_etdff_3/magic_inv_1/Y magic_etdff_2/magic_dff_1/magic_nand_2/Y 4.25e-20
C137 S0 VDD 0.375431f
C138 magic_etdff_0/magic_inv_1/X magic_etdff_0/D 0.027479f
C139 S0 magic_etdff_1/magic_dff_1/D 0.020262f
C140 S3 S1 0.017244f
C141 magic_etdff_2/magic_dff_1/D S1 0.0163f
C142 S1 magic_etdff_1/D 2.325321f
C143 S2 magic_etdff_3/magic_dff_1/D 0.047908f
C144 magic_etdff_3/D magic_etdff_3/magic_dff_1/magic_nand_1/a_100_n230# 0.005219f
C145 S3 VDD 0.008632f
C146 magic_etdff_1/D VDD 0.304704f
C147 magic_etdff_3/magic_dff_0/notQ S1 7.31e-19
C148 magic_etdff_1/magic_dff_1/D magic_etdff_1/D 5.21e-19
C149 magic_etdff_2/magic_dff_1/magic_nand_3/Y magic_etdff_0/magic_dff_1/magic_nand_2/Y 2.01e-20
C150 magic_etdff_3/magic_inv_1/X S1 0.023214f
C151 magic_etdff_3/magic_inv_1/X magic_etdff_2/magic_dff_1/magic_nand_2/Y 0.004704f
C152 magic_etdff_3/magic_inv_1/X VSS 3.119755f
C153 magic_etdff_3/magic_dff_1/D VSS 2.55962f
C154 magic_etdff_3/magic_dff_1/magic_nand_3/Y VSS 0.625399f
C155 magic_etdff_3/magic_dff_1/magic_nand_3/a_100_n230# VSS 0.028228f
C156 magic_etdff_3/magic_dff_1/magic_nand_2/Y VSS 0.662268f
C157 magic_etdff_3/magic_inv_1/Y VSS 3.822167f
C158 magic_etdff_3/magic_dff_1/magic_inv_0/Y VSS 0.535363f
C159 magic_etdff_3/magic_dff_1/magic_nand_2/a_100_n230# VSS 0.028228f
C160 S3 VSS 1.493193f
C161 magic_etdff_3/magic_dff_1/magic_nand_1/a_100_n230# VSS 0.028228f
C162 magic_etdff_3/magic_dff_1/magic_nand_0/a_100_n230# VSS 0.028228f
C163 magic_etdff_3/D VSS 6.593878f
C164 magic_etdff_3/magic_dff_0/magic_nand_3/Y VSS 0.625399f
C165 magic_etdff_3/magic_dff_0/magic_nand_3/a_100_n230# VSS 0.028228f
C166 magic_etdff_3/magic_dff_0/magic_nand_2/Y VSS 0.662029f
C167 magic_etdff_3/magic_dff_0/magic_inv_0/Y VSS 0.53536f
C168 magic_etdff_3/magic_dff_0/magic_nand_2/a_100_n230# VSS 0.028228f
C169 magic_etdff_3/magic_dff_0/magic_nand_1/a_100_n230# VSS 0.028228f
C170 magic_etdff_3/magic_dff_0/notQ VSS 1.07631f
C171 magic_etdff_3/magic_dff_0/magic_nand_0/a_100_n230# VSS 0.028228f
C172 magic_etdff_2/magic_inv_1/X VSS 3.130025f
C173 magic_etdff_2/magic_dff_1/D VSS 2.561133f
C174 magic_etdff_2/magic_dff_1/magic_nand_3/Y VSS 0.627189f
C175 magic_etdff_2/magic_dff_1/magic_nand_3/a_100_n230# VSS 0.028228f
C176 magic_etdff_2/magic_dff_1/magic_nand_2/Y VSS 0.670286f
C177 magic_etdff_2/magic_inv_1/Y VSS 3.826767f
C178 magic_etdff_2/magic_dff_1/magic_inv_0/Y VSS 0.535363f
C179 magic_etdff_2/magic_dff_1/magic_nand_2/a_100_n230# VSS 0.028228f
C180 S2 VSS 3.543593f
C181 magic_etdff_2/magic_dff_1/magic_nand_1/a_100_n230# VSS 0.030804f
C182 magic_etdff_2/magic_dff_1/magic_nand_0/a_100_n230# VSS 0.028228f
C183 magic_etdff_2/D VSS 6.653334f
C184 magic_etdff_2/magic_dff_0/magic_nand_3/Y VSS 0.626657f
C185 magic_etdff_2/magic_dff_0/magic_nand_3/a_100_n230# VSS 0.028228f
C186 magic_etdff_2/magic_dff_0/magic_nand_2/Y VSS 0.662029f
C187 magic_etdff_2/magic_dff_0/magic_inv_0/Y VSS 0.53536f
C188 magic_etdff_2/magic_dff_0/magic_nand_2/a_100_n230# VSS 0.028228f
C189 magic_etdff_2/magic_dff_0/magic_nand_1/a_100_n230# VSS 0.028228f
C190 magic_etdff_2/magic_dff_0/notQ VSS 1.077229f
C191 magic_etdff_2/magic_dff_0/magic_nand_0/a_100_n230# VSS 0.028228f
C192 magic_etdff_1/magic_inv_1/X VSS 3.117251f
C193 VDD VSS 56.242584f
C194 magic_etdff_1/magic_dff_1/D VSS 2.559354f
C195 magic_etdff_1/magic_dff_1/magic_nand_3/Y VSS 0.625399f
C196 magic_etdff_1/magic_dff_1/magic_nand_3/a_100_n230# VSS 0.028228f
C197 magic_etdff_1/magic_dff_1/magic_nand_2/Y VSS 0.6619f
C198 magic_etdff_1/magic_inv_1/Y VSS 3.796575f
C199 magic_etdff_1/magic_dff_1/magic_inv_0/Y VSS 0.535219f
C200 magic_etdff_1/magic_dff_1/magic_nand_2/a_100_n230# VSS 0.028228f
C201 S1 VSS 2.82905f
C202 magic_etdff_1/magic_dff_1/magic_nand_1/a_100_n230# VSS 0.028228f
C203 magic_etdff_1/D VSS 4.68354f
C204 magic_etdff_1/magic_dff_1/magic_nand_0/a_100_n230# VSS 0.028228f
C205 magic_etdff_1/magic_dff_0/magic_nand_3/Y VSS 0.625399f
C206 magic_etdff_1/magic_dff_0/magic_nand_3/a_100_n230# VSS 0.028228f
C207 magic_etdff_1/magic_dff_0/magic_nand_2/Y VSS 0.6619f
C208 magic_etdff_1/magic_dff_0/magic_inv_0/Y VSS 0.535212f
C209 magic_etdff_1/magic_dff_0/magic_nand_2/a_100_n230# VSS 0.028228f
C210 magic_etdff_1/magic_dff_0/magic_nand_1/a_100_n230# VSS 0.028228f
C211 magic_etdff_1/magic_dff_0/notQ VSS 1.07631f
C212 magic_etdff_1/magic_dff_0/magic_nand_0/a_100_n230# VSS 0.028228f
C213 magic_etdff_0/magic_inv_1/X VSS 3.119415f
C214 clk VSS 0.585955f
C215 magic_etdff_0/magic_dff_1/D VSS 2.559354f
C216 magic_etdff_0/magic_dff_1/magic_nand_3/Y VSS 0.625399f
C217 magic_etdff_0/magic_dff_1/magic_nand_3/a_100_n230# VSS 0.028228f
C218 magic_etdff_0/magic_dff_1/magic_nand_2/Y VSS 0.669589f
C219 magic_etdff_0/magic_inv_1/Y VSS 3.797072f
C220 magic_etdff_0/magic_dff_1/magic_inv_0/Y VSS 0.535219f
C221 magic_etdff_0/magic_dff_1/magic_nand_2/a_100_n230# VSS 0.028228f
C222 S0 VSS 5.25179f
C223 magic_etdff_0/magic_dff_1/magic_nand_1/a_100_n230# VSS 0.030804f
C224 magic_etdff_0/D VSS 5.347218f
C225 magic_etdff_0/magic_dff_1/magic_nand_0/a_100_n230# VSS 0.028228f
C226 magic_etdff_0/magic_dff_0/magic_nand_3/Y VSS 0.625399f
C227 magic_etdff_0/magic_dff_0/magic_nand_3/a_100_n230# VSS 0.028228f
C228 magic_etdff_0/magic_dff_0/magic_nand_2/Y VSS 0.6619f
C229 magic_etdff_0/magic_dff_0/magic_inv_0/Y VSS 0.535215f
C230 magic_etdff_0/magic_dff_0/magic_nand_2/a_100_n230# VSS 0.028228f
C231 magic_etdff_0/magic_dff_0/magic_nand_1/a_100_n230# VSS 0.028228f
C232 magic_etdff_0/magic_dff_0/notQ VSS 1.07631f
C233 magic_etdff_0/magic_dff_0/magic_nand_0/a_100_n230# VSS 0.028228f
.ends

.subckt pwm clk S0 S1 S2 S3 PWM VDD VSS
Xmagic_nand_0 magic_nand_0/A magic_nand_0/B magic_nand_1/A VDD VSS magic_nand_0/a_100_n230#
+ magic_nand
Xmagic_nand_1 magic_nand_1/A magic_dff_0/Q magic_nand_1/Y VDD VSS magic_nand_1/a_100_n230#
+ magic_nand
Xmagic_dff_0 magic_comp_0/Y magic_dff_0/Q magic_dff_0/magic_nand_2/Y magic_dff_0/magic_nand_3/Y
+ magic_dff_0/notQ magic_dff_0/magic_nand_1/a_100_n230# magic_dff_0/magic_nand_2/a_100_n230#
+ magic_dff_0/magic_inv_0/Y clk VDD VSS magic_dff
Xmagic_comp_0 magic_comp_0/A0 magic_comp_0/A1 magic_comp_0/Y magic_comp_0/magic_and_1/magic_inv_0/X
+ magic_comp_0/magic_and_1/B magic_comp_0/magic_xnor_1/magic_inv_1/Y magic_comp_0/magic_xnor_1/magic_inv_0/Y
+ magic_comp_0/magic_xnor_0/magic_nand_2/Y magic_comp_0/magic_xnor_2/magic_nand_1/Y
+ magic_comp_0/magic_and_2/magic_inv_0/X magic_comp_0/magic_xnor_2/magic_inv_0/Y magic_comp_0/magic_xnor_2/magic_inv_1/Y
+ magic_comp_0/magic_xnor_3/magic_nand_1/Y magic_nand_0/A magic_comp_0/magic_xnor_1/magic_nand_2/Y
+ magic_comp_0/magic_and_0/B magic_comp_0/magic_xnor_3/magic_nand_0/a_100_n230# S0
+ magic_comp_0/magic_xnor_3/magic_nand_2/Y magic_comp_0/magic_xnor_3/magic_nand_1/a_100_n230#
+ magic_comp_0/magic_and_2/B magic_comp_0/magic_xnor_3/magic_inv_1/Y S3 magic_comp_0/magic_and_1/A
+ magic_comp_0/magic_xnor_0/magic_nand_1/Y magic_comp_0/magic_xnor_3/magic_inv_0/Y
+ magic_comp_0/magic_xnor_2/magic_nand_2/Y magic_comp_0/magic_and_0/magic_inv_0/X
+ magic_comp_0/magic_and_0/A magic_comp_0/magic_xnor_0/magic_inv_1/Y magic_comp_0/magic_xnor_0/magic_inv_0/Y
+ VDD S1 magic_comp_0/A2 magic_comp_0/magic_and_2/A magic_comp_0/magic_xnor_1/magic_nand_1/Y
+ VSS S2 magic_comp
Xmagic_etdff_0 clk magic_etdff_0/magic_dff_1/magic_nand_1/a_100_n230# magic_etdff_0/magic_dff_0/magic_nand_3/Y
+ magic_etdff_0/magic_dff_1/magic_nand_2/a_100_n230# magic_etdff_0/magic_dff_0/magic_inv_0/Y
+ magic_etdff_0/magic_dff_1/magic_nand_3/Y magic_nand_0/B magic_etdff_0/magic_inv_1/Y
+ magic_etdff_0/magic_dff_1/magic_inv_0/Y magic_etdff_0/magic_dff_0/magic_nand_2/Y
+ magic_etdff_0/magic_dff_1/D magic_etdff_0/magic_inv_1/X magic_etdff_0/magic_dff_0/notQ
+ magic_nand_0/A magic_etdff_0/magic_dff_1/magic_nand_2/Y VDD magic_etdff_0/Q VSS
+ magic_etdff
Xmagic_etdff_1 magic_nand_1/Y magic_etdff_1/magic_dff_1/magic_nand_1/a_100_n230# magic_etdff_1/magic_dff_0/magic_nand_3/Y
+ magic_etdff_1/magic_dff_1/magic_nand_2/a_100_n230# magic_etdff_1/magic_dff_0/magic_inv_0/Y
+ magic_etdff_1/magic_dff_1/magic_nand_3/Y magic_etdff_1/D magic_etdff_1/magic_inv_1/Y
+ magic_etdff_1/magic_dff_1/magic_inv_0/Y magic_etdff_1/magic_dff_0/magic_nand_2/Y
+ magic_etdff_1/magic_dff_1/D magic_etdff_1/magic_inv_1/X magic_etdff_1/magic_dff_0/notQ
+ magic_etdff_1/D magic_etdff_1/magic_dff_1/magic_nand_2/Y VDD PWM VSS magic_etdff
Xmagic_counter_0 clk magic_comp_0/A0 magic_comp_0/A1 magic_comp_0/A2 magic_nand_0/A
+ magic_counter_0/magic_etdff_1/magic_dff_1/D magic_counter_0/magic_etdff_0/magic_dff_1/magic_nand_3/Y
+ magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_2/Y magic_counter_0/magic_etdff_2/magic_dff_0/notQ
+ magic_counter_0/magic_etdff_1/magic_inv_1/Y magic_counter_0/magic_etdff_1/magic_dff_1/magic_nand_3/Y
+ magic_counter_0/magic_etdff_2/magic_dff_0/magic_inv_0/Y magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_1/a_100_n230#
+ magic_counter_0/magic_etdff_2/magic_dff_1/D magic_counter_0/magic_etdff_1/magic_inv_1/X
+ magic_counter_0/magic_etdff_3/magic_dff_0/magic_inv_0/Y magic_counter_0/magic_etdff_1/magic_dff_0/notQ
+ magic_counter_0/magic_etdff_2/magic_dff_1/magic_inv_0/Y magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_3/Y
+ magic_counter_0/magic_etdff_2/magic_dff_0/magic_nand_2/Y magic_counter_0/magic_etdff_0/D
+ magic_counter_0/magic_etdff_0/magic_inv_1/Y magic_counter_0/magic_etdff_0/magic_dff_1/D
+ magic_counter_0/magic_etdff_0/magic_inv_1/X magic_counter_0/magic_etdff_3/magic_dff_0/notQ
+ magic_counter_0/magic_etdff_2/D magic_counter_0/magic_etdff_3/magic_dff_1/magic_inv_0/Y
+ magic_counter_0/magic_etdff_0/magic_dff_0/magic_nand_3/Y magic_counter_0/magic_etdff_3/magic_inv_1/X
+ magic_counter_0/magic_etdff_3/magic_inv_1/Y magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_2/Y
+ magic_counter_0/magic_etdff_2/magic_inv_1/X magic_counter_0/magic_etdff_1/D magic_counter_0/magic_etdff_0/magic_dff_0/notQ
+ magic_counter_0/magic_etdff_2/magic_dff_1/magic_nand_2/Y magic_counter_0/magic_etdff_0/magic_dff_0/magic_inv_0/Y
+ magic_counter_0/magic_etdff_3/magic_dff_1/D magic_counter_0/magic_etdff_1/magic_dff_0/magic_nand_3/Y
+ VSS magic_counter_0/magic_etdff_3/D VDD magic_counter_0/magic_etdff_2/magic_inv_1/Y
+ magic_counter
C0 S2 magic_comp_0/magic_and_1/A -0.00392f
C1 S1 S0 0.199423f
C2 magic_etdff_0/magic_dff_0/notQ magic_etdff_0/magic_dff_0/magic_nand_2/Y -2.01e-19
C3 magic_comp_0/magic_and_0/magic_inv_0/X clk 0.034513f
C4 VDD magic_comp_0/magic_and_2/magic_inv_0/X -8.33e-19
C5 VDD magic_dff_0/Q 0.528646f
C6 clk magic_nand_0/B 0.001497f
C7 VDD magic_nand_0/A 0.6057f
C8 magic_etdff_1/magic_dff_1/magic_nand_3/Y magic_etdff_1/D 0.030831f
C9 magic_etdff_1/magic_dff_1/magic_nand_2/Y magic_etdff_1/D 3.74e-20
C10 magic_etdff_1/magic_dff_0/magic_nand_2/Y magic_etdff_1/D 3.74e-20
C11 VDD magic_etdff_1/magic_dff_1/magic_nand_3/Y 4.79e-19
C12 VDD S0 0.002573f
C13 magic_counter_0/magic_etdff_3/D magic_counter_0/magic_etdff_3/magic_inv_1/X -2.22e-34
C14 magic_comp_0/magic_and_0/magic_inv_0/X magic_comp_0/A1 -0.001223f
C15 magic_comp_0/A0 magic_comp_0/magic_xnor_0/magic_nand_1/Y 3.16e-20
C16 magic_etdff_1/magic_dff_0/magic_inv_0/Y magic_nand_1/Y 6.18e-21
C17 magic_comp_0/A0 magic_nand_1/Y 0.575899f
C18 magic_nand_0/B magic_etdff_1/magic_inv_1/X 7.5e-19
C19 magic_comp_0/Y clk 0.41837f
C20 magic_nand_1/Y magic_etdff_1/magic_inv_1/Y 0.100428f
C21 magic_nand_0/A magic_counter_0/magic_etdff_3/magic_inv_1/X 7.14e-19
C22 magic_etdff_1/D magic_nand_1/A 0.001388f
C23 VDD magic_nand_1/a_100_n230# -7.04e-19
C24 clk magic_counter_0/magic_etdff_2/magic_inv_1/Y 0.001371f
C25 S1 clk 0.041558f
C26 magic_comp_0/magic_and_0/magic_inv_0/X magic_comp_0/magic_xnor_1/magic_inv_1/Y -6.54e-19
C27 VDD magic_nand_1/A 0.038267f
C28 S3 magic_counter_0/magic_etdff_2/magic_dff_1/magic_nand_2/Y 0.002756f
C29 magic_etdff_0/magic_dff_1/magic_inv_0/Y magic_etdff_0/magic_dff_0/magic_nand_2/Y -4.14e-19
C30 magic_counter_0/magic_etdff_3/magic_dff_0/notQ magic_comp_0/magic_xnor_3/magic_nand_2/Y 2.83e-20
C31 magic_comp_0/Y magic_dff_0/magic_nand_3/Y 7.19e-19
C32 S2 magic_comp_0/A0 7.25e-19
C33 magic_comp_0/A0 magic_counter_0/magic_etdff_3/magic_dff_1/magic_inv_0/Y 1.38e-19
C34 VDD magic_comp_0/magic_and_1/B -7.85e-19
C35 magic_counter_0/magic_etdff_2/D magic_nand_0/A 1.061227f
C36 magic_comp_0/magic_xnor_2/magic_inv_0/Y magic_comp_0/magic_and_1/magic_inv_0/X -7.57e-19
C37 magic_comp_0/A2 magic_nand_1/Y 1.57e-19
C38 magic_counter_0/magic_etdff_2/magic_inv_1/Y magic_comp_0/A1 1.57e-19
C39 magic_nand_0/B magic_etdff_0/magic_dff_0/magic_nand_2/Y 3.74e-20
C40 magic_etdff_0/Q magic_nand_0/B 0.010221f
C41 S1 magic_comp_0/A1 2.17e-19
C42 VDD clk 1.701662f
C43 magic_counter_0/magic_etdff_3/magic_inv_1/Y S3 0.001513f
C44 S3 magic_counter_0/magic_etdff_3/magic_dff_0/magic_inv_0/Y 0.001074f
C45 magic_dff_0/Q magic_etdff_0/magic_inv_1/X 0.033386f
C46 VDD magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_2/Y 2.99e-19
C47 magic_etdff_1/D magic_comp_0/A1 0.004332f
C48 magic_nand_0/A magic_etdff_0/magic_inv_1/X 0.013108f
C49 magic_etdff_1/D magic_etdff_1/magic_inv_1/X 0.067293f
C50 magic_etdff_0/magic_dff_1/D magic_etdff_0/magic_inv_1/Y -0.049436f
C51 S2 magic_comp_0/A2 2.26e-19
C52 magic_counter_0/magic_etdff_3/magic_dff_1/magic_inv_0/Y magic_comp_0/A2 2.79e-19
C53 VDD magic_dff_0/magic_nand_3/Y 3.35e-20
C54 S3 magic_comp_0/magic_and_2/B -0.001222f
C55 VDD magic_comp_0/A1 1.440218f
C56 magic_comp_0/magic_xnor_1/magic_nand_2/Y clk 0.004896f
C57 VDD magic_etdff_1/magic_inv_1/X 0.006359f
C58 magic_comp_0/magic_xnor_3/magic_inv_0/Y magic_comp_0/Y -1.24e-19
C59 VDD magic_comp_0/magic_xnor_3/magic_nand_2/Y 0.007531f
C60 magic_nand_0/a_100_n230# magic_comp_0/A0 1.35e-19
C61 magic_nand_0/A magic_counter_0/magic_etdff_2/magic_dff_0/notQ 0.001804f
C62 VDD magic_dff_0/notQ -5.15e-19
C63 magic_comp_0/magic_xnor_3/magic_nand_1/Y magic_counter_0/magic_etdff_3/magic_dff_0/notQ 6.69e-22
C64 magic_comp_0/magic_xnor_2/magic_inv_1/Y magic_comp_0/magic_and_1/A -0.001332f
C65 VDD magic_counter_0/magic_etdff_1/magic_dff_1/magic_nand_3/Y 0.004766f
C66 magic_nand_1/a_100_n230# magic_etdff_0/magic_inv_1/X 8.46e-20
C67 VDD magic_comp_0/magic_xnor_1/magic_inv_1/Y -7.6e-19
C68 clk magic_counter_0/magic_etdff_2/D 0.034643f
C69 magic_comp_0/A1 magic_counter_0/magic_etdff_3/magic_inv_1/X 3.03e-19
C70 magic_nand_1/A magic_etdff_0/magic_inv_1/X 0.007345f
C71 magic_counter_0/magic_etdff_3/D magic_nand_1/Y 2.4e-19
C72 magic_comp_0/magic_and_2/B magic_comp_0/magic_xnor_2/magic_inv_0/Y -9.81e-20
C73 VDD magic_etdff_0/Q -3.41e-19
C74 VDD magic_counter_0/magic_etdff_1/magic_dff_0/magic_nand_3/Y 0.004766f
C75 VDD magic_counter_0/magic_etdff_0/magic_inv_1/X 0.007168f
C76 magic_comp_0/magic_and_0/B magic_comp_0/magic_and_0/A -0.001762f
C77 clk magic_comp_0/magic_xnor_1/magic_nand_1/Y 7.46e-20
C78 magic_nand_1/Y magic_dff_0/Q 0.091939f
C79 magic_counter_0/magic_etdff_2/D magic_comp_0/A1 0.042824f
C80 magic_nand_1/Y magic_nand_0/A 0.011639f
C81 VDD magic_comp_0/magic_xnor_0/magic_inv_0/Y -8.48e-19
C82 VDD magic_comp_0/magic_and_1/magic_inv_0/X -8.33e-19
C83 clk magic_etdff_0/magic_inv_1/X 0.007177f
C84 magic_comp_0/A0 magic_comp_0/magic_and_2/A 0.014783f
C85 VDD magic_comp_0/magic_xnor_3/magic_nand_1/Y 0.005259f
C86 magic_comp_0/A2 magic_comp_0/magic_and_1/A -3.19e-19
C87 magic_etdff_0/magic_dff_0/notQ magic_nand_0/B 0.020783f
C88 magic_comp_0/A0 magic_counter_0/magic_etdff_3/magic_dff_1/D 2.97e-19
C89 S2 magic_nand_0/A 1.52e-19
C90 magic_counter_0/magic_etdff_3/magic_dff_1/magic_inv_0/Y magic_nand_0/A 4.54e-19
C91 magic_nand_1/Y magic_nand_1/a_100_n230# -0.013335f
C92 magic_dff_0/notQ magic_etdff_0/magic_inv_1/X 8.86e-21
C93 magic_comp_0/magic_xnor_3/magic_nand_1/Y magic_counter_0/magic_etdff_3/magic_inv_1/X 7.33e-20
C94 magic_comp_0/magic_and_0/magic_inv_0/X magic_comp_0/magic_xnor_1/magic_inv_0/Y -7.57e-19
C95 magic_nand_1/Y magic_nand_1/A 0.033867f
C96 magic_comp_0/A0 magic_etdff_1/magic_inv_1/Y 2.12e-19
C97 VDD magic_counter_0/magic_etdff_3/magic_inv_1/Y 1.38e-19
C98 VDD magic_counter_0/magic_etdff_3/magic_dff_0/magic_inv_0/Y 9.95e-19
C99 magic_counter_0/magic_etdff_3/magic_dff_1/D magic_comp_0/A2 5.7e-19
C100 VDD magic_counter_0/magic_etdff_1/magic_inv_1/Y 0.004482f
C101 clk magic_comp_0/magic_xnor_0/magic_nand_1/Y 7.46e-20
C102 VDD magic_comp_0/magic_and_2/B -7.85e-19
C103 S3 magic_counter_0/magic_etdff_2/magic_inv_1/Y 0.002156f
C104 magic_etdff_0/magic_dff_0/magic_nand_3/Y magic_nand_0/B 0.030353f
C105 VDD magic_counter_0/magic_etdff_1/magic_dff_1/D 0.004724f
C106 magic_comp_0/A0 magic_comp_0/A2 0.037185f
C107 S2 magic_comp_0/magic_and_1/B -0.001222f
C108 VDD magic_comp_0/magic_xnor_3/magic_nand_1/a_100_n230# 7.56e-19
C109 magic_comp_0/A2 magic_etdff_1/magic_inv_1/Y 6.09e-20
C110 VDD magic_etdff_0/magic_dff_0/notQ -3.34e-19
C111 VDD magic_counter_0/magic_etdff_1/magic_dff_0/notQ 0.001384f
C112 magic_nand_1/Y magic_etdff_1/magic_inv_1/X 0.018777f
C113 S2 clk 0.041687f
C114 magic_counter_0/magic_etdff_3/magic_dff_1/magic_inv_0/Y clk 9.19e-20
C115 magic_etdff_0/magic_inv_1/Y magic_dff_0/Q 0.61873f
C116 VDD S3 0.003644f
C117 magic_comp_0/A0 magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_2/Y 3.28e-19
C118 VDD magic_comp_0/magic_xnor_0/magic_inv_1/Y -7.6e-19
C119 VDD magic_comp_0/magic_xnor_1/magic_inv_0/Y -8.48e-19
C120 S2 magic_comp_0/A1 3.71e-19
C121 magic_counter_0/magic_etdff_3/magic_dff_1/magic_inv_0/Y magic_comp_0/A1 1.9e-19
C122 magic_etdff_0/magic_dff_1/D magic_dff_0/Q 0.315289f
C123 magic_comp_0/magic_and_2/A magic_comp_0/magic_and_2/magic_inv_0/X -0.001846f
C124 magic_comp_0/magic_and_2/A magic_comp_0/magic_xnor_3/magic_inv_1/Y -0.001332f
C125 magic_comp_0/magic_and_0/magic_inv_0/X S1 -2.93e-19
C126 magic_counter_0/magic_etdff_3/D magic_counter_0/magic_etdff_3/magic_dff_1/D -2.22e-34
C127 magic_nand_0/A magic_comp_0/magic_and_2/A -3.19e-19
C128 S3 magic_counter_0/magic_etdff_3/magic_inv_1/X 0.004866f
C129 VDD magic_comp_0/magic_xnor_2/magic_inv_0/Y -8.48e-19
C130 clk magic_comp_0/magic_and_0/A 0.285313f
C131 magic_counter_0/magic_etdff_3/magic_dff_1/D magic_nand_0/A 8.54e-19
C132 magic_comp_0/A2 magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_2/Y 6.14e-19
C133 magic_comp_0/A0 magic_counter_0/magic_etdff_3/D 2.83e-19
C134 magic_etdff_0/magic_dff_1/magic_nand_3/Y magic_dff_0/Q 2.5e-19
C135 VDD magic_comp_0/magic_and_0/magic_inv_0/X -8.33e-19
C136 magic_comp_0/magic_and_1/A magic_comp_0/magic_and_1/B -0.001762f
C137 S3 magic_counter_0/magic_etdff_2/D 0.003523f
C138 VDD magic_nand_0/B 0.677177f
C139 magic_comp_0/A0 magic_dff_0/Q 0.003283f
C140 magic_etdff_1/magic_dff_0/magic_inv_0/Y magic_dff_0/Q 3.35e-20
C141 magic_counter_0/magic_etdff_2/magic_dff_1/D magic_nand_0/A 0.016817f
C142 magic_comp_0/A1 magic_comp_0/magic_and_0/A -3.19e-19
C143 magic_dff_0/Q magic_etdff_1/magic_inv_1/Y 0.001945f
C144 magic_comp_0/A0 magic_nand_0/A 1.254507f
C145 clk magic_comp_0/magic_and_1/A 0.293384f
C146 S2 magic_comp_0/magic_and_1/magic_inv_0/X -2.93e-19
C147 magic_comp_0/A0 S0 2.24e-19
C148 VDD magic_comp_0/magic_xnor_3/magic_nand_0/a_100_n230# 7.1e-19
C149 magic_counter_0/magic_etdff_3/D magic_comp_0/A2 7.35e-19
C150 VDD magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_1/a_100_n230# 0.001897f
C151 magic_comp_0/magic_xnor_2/magic_nand_2/Y clk 0.004896f
C152 VDD magic_comp_0/Y 0.011776f
C153 magic_comp_0/magic_xnor_1/magic_inv_1/Y magic_comp_0/magic_and_0/A -0.001332f
C154 clk magic_comp_0/magic_and_2/A 0.342328f
C155 magic_comp_0/A2 magic_nand_0/A 4.339907f
C156 magic_comp_0/magic_xnor_2/magic_inv_1/Y magic_comp_0/magic_and_1/B -0.001122f
C157 VDD S1 7.67e-19
C158 magic_dff_0/notQ magic_etdff_0/magic_inv_1/Y 1.07e-20
C159 magic_nand_0/A magic_counter_0/magic_etdff_2/magic_dff_0/magic_inv_0/Y 0.007393f
C160 magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_2/Y magic_comp_0/magic_and_2/A 2.66e-20
C161 magic_comp_0/A0 magic_nand_1/A 0.005621f
C162 magic_etdff_1/magic_dff_0/magic_inv_0/Y magic_nand_1/A 2.25e-19
C163 magic_counter_0/magic_etdff_3/magic_dff_1/D clk 8.69e-20
C164 magic_etdff_1/magic_inv_1/Y magic_nand_1/A 2.31e-19
C165 magic_comp_0/A2 S0 9.91e-20
C166 magic_comp_0/magic_xnor_2/magic_inv_1/Y clk 0.032672f
C167 VDD magic_etdff_1/D 0.975031f
C168 magic_dff_0/magic_nand_3/Y magic_comp_0/magic_and_2/A 0.001146f
C169 magic_comp_0/magic_and_0/magic_inv_0/X magic_comp_0/magic_xnor_1/magic_nand_1/Y -3.43e-20
C170 magic_comp_0/Y magic_dff_0/magic_inv_0/Y 0.001473f
C171 magic_counter_0/magic_etdff_2/magic_dff_0/magic_nand_2/Y magic_nand_0/A 0.007076f
C172 magic_comp_0/A0 clk 0.56752f
C173 magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_2/Y magic_nand_0/A 0.00258f
C174 magic_etdff_0/magic_inv_1/Y magic_etdff_0/magic_dff_0/magic_nand_2/Y -0.011355f
C175 magic_counter_0/magic_etdff_3/magic_dff_1/D magic_comp_0/A1 3.87e-19
C176 magic_etdff_1/D magic_etdff_1/magic_dff_0/notQ 0.020796f
C177 magic_nand_0/B magic_etdff_0/magic_inv_1/X 0.052326f
C178 magic_comp_0/A0 magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_2/Y 1.11e-19
C179 VDD magic_etdff_1/magic_dff_0/notQ 2.66e-20
C180 magic_comp_0/magic_and_1/A magic_comp_0/magic_and_1/magic_inv_0/X -0.001846f
C181 magic_comp_0/A0 magic_dff_0/magic_nand_3/Y 2.11e-20
C182 magic_comp_0/A0 magic_comp_0/A1 5.97106f
C183 magic_comp_0/A0 magic_etdff_1/magic_inv_1/X 0.016848f
C184 magic_etdff_0/magic_dff_1/D magic_etdff_0/magic_dff_0/magic_nand_2/Y -1.04e-20
C185 VDD magic_counter_0/magic_etdff_3/magic_inv_1/X 4.07e-19
C186 magic_comp_0/A0 magic_comp_0/magic_xnor_3/magic_nand_2/Y 0.004578f
C187 magic_comp_0/magic_xnor_3/magic_inv_0/Y magic_comp_0/magic_and_2/A -0.00139f
C188 magic_dff_0/notQ magic_comp_0/A0 2.11e-20
C189 magic_comp_0/A2 clk 0.01474f
C190 magic_counter_0/magic_etdff_3/D magic_nand_0/A 2.1938f
C191 S2 S3 0.199423f
C192 clk magic_counter_0/magic_etdff_2/magic_dff_0/magic_inv_0/Y 4.14e-20
C193 magic_comp_0/magic_and_2/magic_inv_0/X magic_comp_0/magic_xnor_3/magic_inv_1/Y -6.54e-19
C194 VDD magic_counter_0/magic_etdff_1/D 0.007441f
C195 magic_comp_0/magic_and_0/B clk 0.074404f
C196 magic_comp_0/A2 magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_2/Y 2.39e-19
C197 magic_nand_0/A magic_comp_0/magic_and_2/magic_inv_0/X -0.001223f
C198 VDD magic_counter_0/magic_etdff_2/D 8.7e-20
C199 magic_nand_0/A magic_dff_0/Q 0.013967f
C200 magic_comp_0/A2 magic_comp_0/A1 4.993299f
C201 magic_comp_0/A2 magic_etdff_1/magic_inv_1/X 4.27e-20
C202 magic_comp_0/magic_xnor_2/magic_inv_1/Y magic_comp_0/magic_and_1/magic_inv_0/X -6.54e-19
C203 magic_comp_0/A2 magic_comp_0/magic_xnor_3/magic_nand_2/Y 1.52e-19
C204 magic_comp_0/magic_xnor_3/magic_nand_1/Y magic_counter_0/magic_etdff_3/magic_dff_1/D 0.00147f
C205 magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_2/Y clk 7.12e-20
C206 magic_nand_0/A S0 7.31e-20
C207 magic_nand_1/Y magic_nand_0/B 0.010394f
C208 VDD magic_counter_0/magic_etdff_0/magic_dff_1/D 0.004724f
C209 VDD magic_etdff_0/magic_inv_1/X 0.005572f
C210 VDD magic_counter_0/magic_etdff_0/magic_dff_1/magic_nand_3/Y 0.004766f
C211 clk magic_counter_0/magic_etdff_0/magic_dff_0/magic_inv_0/Y 4.14e-20
C212 magic_comp_0/magic_xnor_3/magic_nand_1/Y magic_comp_0/A0 0.018694f
C213 magic_counter_0/magic_etdff_0/magic_inv_1/Y clk 0.001371f
C214 magic_nand_1/a_100_n230# magic_dff_0/Q 0.038264f
C215 magic_etdff_0/magic_dff_1/magic_nand_2/Y magic_dff_0/Q 1.52e-19
C216 VDD magic_counter_0/magic_etdff_0/magic_dff_0/notQ 0.001384f
C217 magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_2/Y magic_comp_0/A1 4.37e-19
C218 magic_dff_0/Q magic_nand_1/A 0.061152f
C219 magic_comp_0/magic_and_0/B magic_comp_0/magic_xnor_1/magic_inv_1/Y -0.001122f
C220 magic_nand_0/A magic_nand_1/A 1.47e-19
C221 magic_etdff_0/magic_dff_0/notQ magic_etdff_0/magic_inv_1/Y -0.018386f
C222 magic_counter_0/magic_etdff_0/D clk 0.035695f
C223 magic_comp_0/magic_xnor_1/magic_inv_0/Y magic_comp_0/magic_and_0/A -0.00139f
C224 magic_counter_0/magic_etdff_3/D clk 7.51e-20
C225 magic_comp_0/A0 magic_counter_0/magic_etdff_2/magic_dff_1/magic_nand_2/Y 1.11e-19
C226 magic_comp_0/magic_and_2/B magic_comp_0/magic_and_2/A -0.001762f
C227 magic_comp_0/A2 magic_comp_0/magic_and_1/magic_inv_0/X -0.001223f
C228 clk magic_comp_0/magic_and_2/magic_inv_0/X 0.034831f
C229 clk magic_comp_0/magic_xnor_3/magic_inv_1/Y 0.044539f
C230 clk magic_dff_0/Q 0.001499f
C231 magic_comp_0/magic_xnor_3/magic_nand_1/Y magic_comp_0/A2 1.89e-19
C232 clk magic_nand_0/A 0.40967f
C233 magic_etdff_0/magic_dff_0/notQ magic_etdff_0/magic_dff_1/D -9.13e-19
C234 magic_counter_0/magic_etdff_3/D magic_comp_0/A1 3.63e-19
C235 magic_counter_0/magic_etdff_3/D magic_etdff_1/magic_inv_1/X 3.36e-19
C236 magic_nand_1/Y magic_etdff_1/D 0.139652f
C237 magic_counter_0/magic_etdff_3/magic_inv_1/Y magic_comp_0/A0 1.38e-19
C238 magic_comp_0/A0 magic_counter_0/magic_etdff_3/magic_dff_0/magic_inv_0/Y 1.38e-19
C239 magic_nand_1/a_100_n230# magic_nand_1/A 3.25e-20
C240 magic_counter_0/magic_etdff_3/D magic_comp_0/magic_xnor_3/magic_nand_2/Y 8.24e-20
C241 magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_2/Y magic_nand_0/A 5.06e-19
C242 magic_comp_0/magic_xnor_2/magic_inv_1/Y magic_comp_0/magic_and_2/B -7.65e-20
C243 clk S0 0.062858f
C244 magic_comp_0/magic_and_0/magic_inv_0/X magic_comp_0/magic_and_0/A -0.001846f
C245 magic_dff_0/magic_nand_3/Y magic_dff_0/Q 4.19e-20
C246 S3 magic_comp_0/magic_and_2/A -0.00392f
C247 VDD magic_nand_1/Y 0.28258f
C248 magic_comp_0/A2 magic_counter_0/magic_etdff_2/magic_dff_1/magic_nand_2/Y 2.39e-19
C249 S2 S1 0.199423f
C250 magic_dff_0/Q magic_etdff_1/magic_inv_1/X 1.23e-19
C251 magic_nand_0/a_100_n230# magic_nand_0/B -1.78e-33
C252 magic_nand_0/A magic_comp_0/A1 0.17683f
C253 magic_nand_0/A magic_etdff_1/magic_inv_1/X 5.53e-19
C254 magic_nand_0/A magic_comp_0/magic_xnor_3/magic_nand_2/Y 1.08e-19
C255 magic_comp_0/magic_xnor_2/magic_inv_0/Y magic_comp_0/magic_and_1/A -0.00139f
C256 magic_dff_0/notQ magic_dff_0/Q 0.003567f
C257 magic_etdff_0/magic_dff_0/magic_nand_3/Y magic_etdff_0/magic_inv_1/Y -1.59e-19
C258 S0 magic_comp_0/A1 1.42e-19
C259 magic_counter_0/magic_etdff_3/magic_inv_1/Y magic_comp_0/A2 2.82e-19
C260 magic_comp_0/A2 magic_counter_0/magic_etdff_3/magic_dff_0/magic_inv_0/Y 2.79e-19
C261 VDD S2 7.67e-19
C262 VDD magic_counter_0/magic_etdff_3/magic_dff_1/magic_inv_0/Y 1.39e-19
C263 magic_etdff_0/magic_inv_1/Y magic_nand_0/B 0.045194f
C264 clk magic_comp_0/magic_and_1/B 0.033079f
C265 magic_comp_0/A0 S3 1.348609f
C266 magic_dff_0/Q magic_etdff_0/magic_dff_0/magic_nand_2/Y 0.029105f
C267 magic_comp_0/magic_xnor_3/magic_inv_0/Y magic_comp_0/magic_and_2/magic_inv_0/X -7.57e-19
C268 S1 magic_comp_0/magic_and_0/A -0.00392f
C269 magic_comp_0/magic_xnor_3/magic_nand_1/Y magic_counter_0/magic_etdff_3/D 1.08e-19
C270 magic_etdff_1/magic_inv_1/X magic_nand_1/A 3.36e-19
C271 magic_counter_0/magic_etdff_2/magic_dff_1/magic_inv_0/Y magic_nand_0/A 0.007393f
C272 magic_etdff_0/magic_dff_1/D magic_nand_0/B 0.034328f
C273 magic_comp_0/magic_xnor_3/magic_nand_1/Y magic_comp_0/magic_and_2/magic_inv_0/X -3.43e-20
C274 magic_nand_0/A magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_3/Y 1.26e-19
C275 magic_comp_0/magic_xnor_3/magic_nand_1/Y magic_nand_0/A 1.38e-19
C276 VDD magic_comp_0/magic_and_0/A -1.27e-19
C277 magic_dff_0/magic_nand_3/Y clk 0.002002f
C278 S3 magic_comp_0/A2 0.027569f
C279 magic_etdff_1/magic_dff_1/D magic_etdff_1/D 0.035054f
C280 clk magic_comp_0/A1 0.033104f
C281 VDD magic_nand_0/a_100_n230# 0.003967f
C282 clk magic_comp_0/magic_xnor_3/magic_nand_2/Y 0.021149f
C283 VDD magic_etdff_1/magic_dff_1/D 4.57e-19
C284 magic_dff_0/notQ clk 2.28e-19
C285 magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_2/Y magic_comp_0/A1 1.57e-19
C286 magic_etdff_0/magic_dff_1/magic_nand_3/Y magic_nand_0/B 0.030353f
C287 magic_comp_0/magic_xnor_1/magic_inv_1/Y magic_comp_0/magic_and_1/B -7.65e-20
C288 magic_comp_0/Y magic_comp_0/magic_and_2/A 0.231885f
C289 clk magic_comp_0/magic_xnor_0/magic_nand_2/Y 0.007048f
C290 magic_nand_0/A magic_counter_0/magic_etdff_2/magic_dff_1/magic_nand_2/Y 4.73e-19
C291 magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_2/Y magic_comp_0/magic_xnor_3/magic_nand_2/Y 0.001256f
C292 magic_nand_0/A magic_counter_0/magic_etdff_2/magic_inv_1/X 0.016149f
C293 magic_comp_0/A0 magic_nand_0/B 0.00795f
C294 magic_nand_0/B magic_etdff_1/magic_inv_1/Y 1.87e-19
C295 magic_comp_0/A1 magic_etdff_1/magic_inv_1/X 7.33e-19
C296 VDD magic_comp_0/magic_and_1/A -1.27e-19
C297 magic_comp_0/magic_xnor_1/magic_inv_1/Y clk 0.032672f
C298 VDD magic_etdff_0/magic_inv_1/Y -0.022882f
C299 magic_comp_0/A1 magic_comp_0/magic_xnor_3/magic_nand_2/Y 2.3e-19
C300 magic_counter_0/magic_etdff_3/magic_inv_1/Y magic_nand_0/A 5.24e-19
C301 magic_counter_0/magic_etdff_3/magic_dff_0/magic_inv_0/Y magic_nand_0/A 4.54e-19
C302 magic_comp_0/magic_xnor_2/magic_nand_1/Y clk 7.46e-20
C303 magic_comp_0/magic_xnor_3/magic_inv_0/Y clk 0.021438f
C304 magic_counter_0/magic_etdff_0/magic_inv_1/X clk 0.029804f
C305 magic_comp_0/A0 magic_comp_0/Y 2.11e-20
C306 VDD magic_etdff_0/magic_dff_1/D -1.29e-19
C307 magic_comp_0/magic_and_2/B magic_comp_0/magic_xnor_3/magic_inv_1/Y -0.001122f
C308 VDD magic_comp_0/magic_and_2/A 0.025334f
C309 clk magic_comp_0/magic_and_1/magic_inv_0/X 0.034513f
C310 clk magic_comp_0/magic_xnor_0/magic_inv_0/Y 0.02115f
C311 magic_comp_0/magic_xnor_3/magic_nand_1/Y clk 5.14e-19
C312 magic_etdff_1/D magic_etdff_1/magic_dff_0/magic_nand_3/Y 0.03094f
C313 magic_comp_0/A0 magic_counter_0/magic_etdff_2/magic_inv_1/Y 1.11e-19
C314 magic_comp_0/A0 S1 3.69e-19
C315 magic_etdff_0/magic_dff_0/notQ magic_dff_0/Q 0.126658f
C316 S3 magic_counter_0/magic_etdff_3/D 0.005527f
C317 VDD magic_counter_0/magic_etdff_3/magic_dff_1/D 9.51e-19
C318 magic_comp_0/magic_xnor_3/magic_nand_1/Y magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_2/Y 4.45e-21
C319 VDD magic_etdff_1/magic_dff_0/magic_nand_3/Y 4.79e-19
C320 VDD magic_comp_0/magic_xnor_2/magic_inv_1/Y -7.6e-19
C321 S3 magic_comp_0/magic_and_2/magic_inv_0/X -2.93e-19
C322 magic_comp_0/A0 magic_etdff_1/D 0.051668f
C323 magic_nand_0/a_100_n230# magic_etdff_0/magic_inv_1/X 0.001946f
C324 clk magic_counter_0/magic_etdff_2/magic_inv_1/X 0.03018f
C325 magic_comp_0/magic_xnor_3/magic_nand_1/Y magic_comp_0/A1 2.76e-19
C326 magic_etdff_1/D magic_etdff_1/magic_inv_1/Y 0.045519f
C327 S3 magic_nand_0/A 0.010158f
C328 VDD magic_etdff_1/magic_dff_0/magic_inv_0/Y 4e-19
C329 VDD magic_comp_0/A0 1.976874f
C330 VDD magic_etdff_1/magic_inv_1/Y 0.007458f
C331 magic_comp_0/A2 magic_counter_0/magic_etdff_2/magic_inv_1/Y 2.39e-19
C332 VDD magic_counter_0/magic_etdff_1/magic_inv_1/X 0.007168f
C333 S1 magic_comp_0/A2 1.47e-19
C334 magic_comp_0/A1 magic_counter_0/magic_etdff_2/magic_dff_1/magic_nand_2/Y 1.57e-19
C335 magic_counter_0/magic_etdff_3/magic_inv_1/Y clk 1.03e-19
C336 magic_comp_0/magic_and_0/B S1 -0.001222f
C337 magic_comp_0/magic_xnor_2/magic_nand_1/Y magic_comp_0/magic_and_1/magic_inv_0/X -3.43e-20
C338 magic_comp_0/A0 magic_counter_0/magic_etdff_3/magic_inv_1/X 2.27e-19
C339 magic_etdff_0/magic_dff_1/magic_inv_0/Y magic_dff_0/Q 0.001199f
C340 magic_etdff_0/magic_dff_0/magic_nand_3/Y magic_dff_0/Q 0.034448f
C341 magic_comp_0/magic_and_2/B clk 0.033079f
C342 VDD magic_comp_0/A2 0.604789f
C343 magic_etdff_0/magic_dff_0/magic_nand_3/Y magic_nand_0/A 1.11e-19
C344 PWM magic_etdff_1/D 0.010894f
C345 magic_counter_0/magic_etdff_3/magic_inv_1/Y magic_comp_0/A1 1.91e-19
C346 magic_counter_0/magic_etdff_3/magic_dff_0/magic_inv_0/Y magic_comp_0/A1 1.9e-19
C347 magic_counter_0/magic_etdff_3/magic_inv_1/Y magic_comp_0/magic_xnor_3/magic_nand_2/Y 6.35e-20
C348 VDD magic_comp_0/magic_and_0/B -7.85e-19
C349 magic_comp_0/A0 magic_counter_0/magic_etdff_1/D 9.81e-20
C350 magic_nand_0/B magic_dff_0/Q 0.230921f
C351 VDD PWM 0.004233f
C352 magic_comp_0/A0 magic_counter_0/magic_etdff_2/D 0.022896f
C353 magic_nand_0/B magic_nand_0/A 0.073251f
C354 S3 clk 0.053093f
C355 magic_comp_0/magic_xnor_1/magic_inv_0/Y magic_comp_0/magic_and_1/B -9.81e-20
C356 magic_comp_0/A2 magic_counter_0/magic_etdff_3/magic_inv_1/X 4.73e-19
C357 VDD magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_2/Y 0.005882f
C358 magic_comp_0/magic_xnor_0/magic_inv_1/Y clk 0.046312f
C359 S3 magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_2/Y 2.68e-21
C360 magic_comp_0/Y magic_comp_0/magic_and_2/magic_inv_0/X 0.004948f
C361 magic_comp_0/Y magic_comp_0/magic_xnor_3/magic_inv_1/Y 0.001077f
C362 magic_comp_0/Y magic_dff_0/Q 2.03e-24
C363 clk magic_comp_0/magic_xnor_1/magic_inv_0/Y 0.021133f
C364 magic_comp_0/A0 magic_etdff_0/magic_inv_1/X 0.002963f
C365 magic_comp_0/Y magic_nand_0/A 1.46e-20
C366 VDD magic_counter_0/magic_etdff_0/magic_inv_1/Y 0.004482f
C367 S3 magic_comp_0/A1 0.041703f
C368 magic_comp_0/A2 magic_counter_0/magic_etdff_2/D 0.093921f
C369 magic_etdff_0/magic_dff_1/magic_nand_2/Y magic_nand_0/B 3.74e-20
C370 VDD magic_counter_0/magic_etdff_0/magic_dff_0/magic_nand_3/Y 0.004766f
C371 magic_nand_0/B magic_nand_1/A 0.022405f
C372 magic_nand_0/A magic_counter_0/magic_etdff_2/magic_inv_1/Y 0.036485f
C373 S1 magic_nand_0/A 1.02e-19
C374 magic_etdff_0/magic_dff_0/magic_inv_0/Y magic_dff_0/Q 0.009506f
C375 VDD magic_counter_0/magic_etdff_0/D 0.002827f
C376 clk magic_comp_0/magic_xnor_2/magic_inv_0/Y 0.021133f
C377 magic_counter_0/magic_etdff_3/magic_inv_1/Y magic_comp_0/magic_xnor_3/magic_nand_1/Y 8.55e-20
C378 VDD magic_counter_0/magic_etdff_3/D 0.009302f
C379 magic_counter_0/magic_etdff_3/magic_inv_1/X VSS 3.121172f
C380 magic_counter_0/magic_etdff_3/magic_dff_1/D VSS 2.559354f
C381 magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_3/Y VSS 0.625399f
C382 magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_3/a_100_n230# VSS 0.028228f
C383 magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_2/Y VSS 0.662089f
C384 magic_counter_0/magic_etdff_3/magic_inv_1/Y VSS 3.797556f
C385 magic_counter_0/magic_etdff_3/magic_dff_1/magic_inv_0/Y VSS 0.535219f
C386 magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_2/a_100_n230# VSS 0.028228f
C387 magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_1/a_100_n230# VSS 0.028228f
C388 magic_counter_0/magic_etdff_3/magic_dff_1/magic_nand_0/a_100_n230# VSS 0.028228f
C389 magic_counter_0/magic_etdff_3/D VSS 4.664954f
C390 magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_3/Y VSS 0.625399f
C391 magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_3/a_100_n230# VSS 0.028228f
C392 magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_2/Y VSS 0.6619f
C393 magic_counter_0/magic_etdff_3/magic_dff_0/magic_inv_0/Y VSS 0.535219f
C394 magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_2/a_100_n230# VSS 0.028228f
C395 magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_1/a_100_n230# VSS 0.028228f
C396 magic_counter_0/magic_etdff_3/magic_dff_0/notQ VSS 1.07631f
C397 magic_counter_0/magic_etdff_3/magic_dff_0/magic_nand_0/a_100_n230# VSS 0.028228f
C398 magic_counter_0/magic_etdff_2/magic_inv_1/X VSS 3.121172f
C399 magic_counter_0/magic_etdff_2/magic_dff_1/D VSS 2.559354f
C400 magic_counter_0/magic_etdff_2/magic_dff_1/magic_nand_3/Y VSS 0.625399f
C401 magic_counter_0/magic_etdff_2/magic_dff_1/magic_nand_3/a_100_n230# VSS 0.028228f
C402 magic_counter_0/magic_etdff_2/magic_dff_1/magic_nand_2/Y VSS 0.6619f
C403 magic_counter_0/magic_etdff_2/magic_inv_1/Y VSS 3.797556f
C404 magic_counter_0/magic_etdff_2/magic_dff_1/magic_inv_0/Y VSS 0.535219f
C405 magic_counter_0/magic_etdff_2/magic_dff_1/magic_nand_2/a_100_n230# VSS 0.028228f
C406 magic_comp_0/A2 VSS 6.68854f
C407 magic_counter_0/magic_etdff_2/magic_dff_1/magic_nand_1/a_100_n230# VSS 0.028228f
C408 magic_counter_0/magic_etdff_2/magic_dff_1/magic_nand_0/a_100_n230# VSS 0.028228f
C409 magic_counter_0/magic_etdff_2/D VSS 4.710068f
C410 magic_counter_0/magic_etdff_2/magic_dff_0/magic_nand_3/Y VSS 0.625399f
C411 magic_counter_0/magic_etdff_2/magic_dff_0/magic_nand_3/a_100_n230# VSS 0.028228f
C412 magic_counter_0/magic_etdff_2/magic_dff_0/magic_nand_2/Y VSS 0.6619f
C413 magic_counter_0/magic_etdff_2/magic_dff_0/magic_inv_0/Y VSS 0.535219f
C414 magic_counter_0/magic_etdff_2/magic_dff_0/magic_nand_2/a_100_n230# VSS 0.028228f
C415 magic_counter_0/magic_etdff_2/magic_dff_0/magic_nand_1/a_100_n230# VSS 0.028228f
C416 magic_counter_0/magic_etdff_2/magic_dff_0/notQ VSS 1.07631f
C417 magic_counter_0/magic_etdff_2/magic_dff_0/magic_nand_0/a_100_n230# VSS 0.028228f
C418 magic_counter_0/magic_etdff_1/magic_inv_1/X VSS 3.121172f
C419 VDD VSS 0.121727p
C420 magic_counter_0/magic_etdff_1/magic_dff_1/D VSS 2.559354f
C421 magic_counter_0/magic_etdff_1/magic_dff_1/magic_nand_3/Y VSS 0.625399f
C422 magic_counter_0/magic_etdff_1/magic_dff_1/magic_nand_3/a_100_n230# VSS 0.028228f
C423 magic_counter_0/magic_etdff_1/magic_dff_1/magic_nand_2/Y VSS 0.6619f
C424 magic_counter_0/magic_etdff_1/magic_inv_1/Y VSS 3.797556f
C425 magic_counter_0/magic_etdff_1/magic_dff_1/magic_inv_0/Y VSS 0.535219f
C426 magic_counter_0/magic_etdff_1/magic_dff_1/magic_nand_2/a_100_n230# VSS 0.028228f
C427 magic_comp_0/A1 VSS 5.189204f
C428 magic_counter_0/magic_etdff_1/magic_dff_1/magic_nand_1/a_100_n230# VSS 0.028228f
C429 magic_counter_0/magic_etdff_1/D VSS 3.137679f
C430 magic_counter_0/magic_etdff_1/magic_dff_1/magic_nand_0/a_100_n230# VSS 0.028228f
C431 magic_counter_0/magic_etdff_1/magic_dff_0/magic_nand_3/Y VSS 0.625399f
C432 magic_counter_0/magic_etdff_1/magic_dff_0/magic_nand_3/a_100_n230# VSS 0.028228f
C433 magic_counter_0/magic_etdff_1/magic_dff_0/magic_nand_2/Y VSS 0.6619f
C434 magic_counter_0/magic_etdff_1/magic_dff_0/magic_inv_0/Y VSS 0.535219f
C435 magic_counter_0/magic_etdff_1/magic_dff_0/magic_nand_2/a_100_n230# VSS 0.028228f
C436 magic_counter_0/magic_etdff_1/magic_dff_0/magic_nand_1/a_100_n230# VSS 0.028228f
C437 magic_counter_0/magic_etdff_1/magic_dff_0/notQ VSS 1.07631f
C438 magic_counter_0/magic_etdff_1/magic_dff_0/magic_nand_0/a_100_n230# VSS 0.028228f
C439 magic_counter_0/magic_etdff_0/magic_inv_1/X VSS 3.121172f
C440 magic_counter_0/magic_etdff_0/magic_dff_1/D VSS 2.559354f
C441 magic_counter_0/magic_etdff_0/magic_dff_1/magic_nand_3/Y VSS 0.625399f
C442 magic_counter_0/magic_etdff_0/magic_dff_1/magic_nand_3/a_100_n230# VSS 0.028228f
C443 magic_counter_0/magic_etdff_0/magic_dff_1/magic_nand_2/Y VSS 0.6619f
C444 magic_counter_0/magic_etdff_0/magic_inv_1/Y VSS 3.797556f
C445 magic_counter_0/magic_etdff_0/magic_dff_1/magic_inv_0/Y VSS 0.535219f
C446 magic_counter_0/magic_etdff_0/magic_dff_1/magic_nand_2/a_100_n230# VSS 0.028228f
C447 magic_comp_0/A0 VSS 7.629625f
C448 magic_counter_0/magic_etdff_0/magic_dff_1/magic_nand_1/a_100_n230# VSS 0.028228f
C449 magic_counter_0/magic_etdff_0/D VSS 3.753388f
C450 magic_counter_0/magic_etdff_0/magic_dff_1/magic_nand_0/a_100_n230# VSS 0.028228f
C451 magic_counter_0/magic_etdff_0/magic_dff_0/magic_nand_3/Y VSS 0.625399f
C452 magic_counter_0/magic_etdff_0/magic_dff_0/magic_nand_3/a_100_n230# VSS 0.028228f
C453 magic_counter_0/magic_etdff_0/magic_dff_0/magic_nand_2/Y VSS 0.6619f
C454 magic_counter_0/magic_etdff_0/magic_dff_0/magic_inv_0/Y VSS 0.535219f
C455 magic_counter_0/magic_etdff_0/magic_dff_0/magic_nand_2/a_100_n230# VSS 0.028228f
C456 magic_counter_0/magic_etdff_0/magic_dff_0/magic_nand_1/a_100_n230# VSS 0.028228f
C457 magic_counter_0/magic_etdff_0/magic_dff_0/notQ VSS 1.07631f
C458 magic_counter_0/magic_etdff_0/magic_dff_0/magic_nand_0/a_100_n230# VSS 0.028228f
C459 magic_etdff_1/magic_inv_1/X VSS 3.12185f
C460 magic_nand_1/Y VSS 1.891323f
C461 magic_etdff_1/magic_dff_1/D VSS 2.559354f
C462 magic_etdff_1/magic_dff_1/magic_nand_3/Y VSS 0.625399f
C463 magic_etdff_1/magic_dff_1/magic_nand_3/a_100_n230# VSS 0.028228f
C464 magic_etdff_1/magic_dff_1/magic_nand_2/Y VSS 0.6619f
C465 magic_etdff_1/magic_inv_1/Y VSS 3.807182f
C466 magic_etdff_1/magic_dff_1/magic_inv_0/Y VSS 0.535219f
C467 magic_etdff_1/magic_dff_1/magic_nand_2/a_100_n230# VSS 0.028228f
C468 PWM VSS 1.470301f
C469 magic_etdff_1/magic_dff_1/magic_nand_1/a_100_n230# VSS 0.028228f
C470 magic_etdff_1/magic_dff_1/magic_nand_0/a_100_n230# VSS 0.028228f
C471 magic_etdff_1/D VSS 6.121228f
C472 magic_etdff_1/magic_dff_0/magic_nand_3/Y VSS 0.625399f
C473 magic_etdff_1/magic_dff_0/magic_nand_3/a_100_n230# VSS 0.028228f
C474 magic_etdff_1/magic_dff_0/magic_nand_2/Y VSS 0.6619f
C475 magic_etdff_1/magic_dff_0/magic_inv_0/Y VSS 0.535219f
C476 magic_etdff_1/magic_dff_0/magic_nand_2/a_100_n230# VSS 0.028228f
C477 magic_etdff_1/magic_dff_0/magic_nand_1/a_100_n230# VSS 0.028228f
C478 magic_etdff_1/magic_dff_0/notQ VSS 1.07631f
C479 magic_etdff_1/magic_dff_0/magic_nand_0/a_100_n230# VSS 0.028228f
C480 magic_etdff_0/magic_inv_1/X VSS 3.126472f
C481 magic_etdff_0/magic_dff_1/D VSS 2.559304f
C482 magic_etdff_0/magic_dff_1/magic_nand_3/Y VSS 0.625399f
C483 magic_etdff_0/magic_dff_1/magic_nand_3/a_100_n230# VSS 0.028228f
C484 magic_etdff_0/magic_dff_1/magic_nand_2/Y VSS 0.677795f
C485 magic_etdff_0/magic_inv_1/Y VSS 3.796909f
C486 magic_etdff_0/magic_dff_1/magic_inv_0/Y VSS 0.535219f
C487 magic_etdff_0/magic_dff_1/magic_nand_2/a_100_n230# VSS 0.028228f
C488 magic_etdff_0/Q VSS 1.461477f
C489 magic_etdff_0/magic_dff_1/magic_nand_1/a_100_n230# VSS 0.032543f
C490 magic_nand_0/B VSS 4.263944f
C491 magic_etdff_0/magic_dff_1/magic_nand_0/a_100_n230# VSS 0.028228f
C492 magic_etdff_0/magic_dff_0/magic_nand_3/Y VSS 0.625399f
C493 magic_etdff_0/magic_dff_0/magic_nand_3/a_100_n230# VSS 0.028228f
C494 magic_etdff_0/magic_dff_0/magic_nand_2/Y VSS 0.661866f
C495 magic_etdff_0/magic_dff_0/magic_inv_0/Y VSS 0.535219f
C496 magic_etdff_0/magic_dff_0/magic_nand_2/a_100_n230# VSS 0.028228f
C497 magic_etdff_0/magic_dff_0/magic_nand_1/a_100_n230# VSS 0.028228f
C498 magic_etdff_0/magic_dff_0/notQ VSS 1.07631f
C499 magic_etdff_0/magic_dff_0/magic_nand_0/a_100_n230# VSS 0.028228f
C500 magic_comp_0/magic_and_2/magic_inv_0/X VSS 0.651385f
C501 magic_comp_0/magic_and_2/B VSS 1.00746f
C502 magic_comp_0/magic_and_2/magic_nand_0/a_100_n230# VSS 0.028228f
C503 magic_comp_0/magic_and_1/magic_inv_0/X VSS 0.65138f
C504 magic_comp_0/magic_and_1/B VSS 1.00746f
C505 magic_comp_0/magic_and_1/magic_nand_0/a_100_n230# VSS 0.028228f
C506 magic_comp_0/magic_and_0/magic_inv_0/X VSS 0.65138f
C507 magic_comp_0/magic_and_0/magic_nand_0/a_100_n230# VSS 0.028228f
C508 magic_comp_0/magic_xnor_3/magic_nand_2/Y VSS 0.736068f
C509 magic_comp_0/magic_xnor_3/magic_inv_1/Y VSS 0.876506f
C510 magic_comp_0/magic_xnor_3/magic_inv_0/Y VSS 0.513303f
C511 magic_comp_0/magic_xnor_3/magic_nand_2/a_100_n230# VSS 0.028228f
C512 magic_comp_0/magic_xnor_3/magic_nand_1/Y VSS 0.570384f
C513 magic_nand_0/A VSS 10.197869f
C514 S3 VSS 2.792103f
C515 magic_comp_0/magic_xnor_3/magic_nand_1/a_100_n230# VSS 0.028228f
C516 magic_comp_0/magic_and_2/A VSS 1.741955f
C517 magic_comp_0/magic_xnor_3/magic_nand_0/a_100_n230# VSS 0.028228f
C518 magic_comp_0/magic_xnor_2/magic_nand_2/Y VSS 0.735869f
C519 magic_comp_0/magic_xnor_2/magic_inv_1/Y VSS 0.876506f
C520 magic_comp_0/magic_xnor_2/magic_inv_0/Y VSS 0.513834f
C521 magic_comp_0/magic_xnor_2/magic_nand_2/a_100_n230# VSS 0.028228f
C522 magic_comp_0/magic_xnor_2/magic_nand_1/Y VSS 0.570102f
C523 S2 VSS 2.433005f
C524 magic_comp_0/magic_xnor_2/magic_nand_1/a_100_n230# VSS 0.028228f
C525 magic_comp_0/magic_and_1/A VSS 1.547636f
C526 magic_comp_0/magic_xnor_2/magic_nand_0/a_100_n230# VSS 0.028228f
C527 magic_comp_0/magic_xnor_1/magic_nand_2/Y VSS 0.735869f
C528 magic_comp_0/magic_xnor_1/magic_inv_1/Y VSS 0.876506f
C529 magic_comp_0/magic_xnor_1/magic_inv_0/Y VSS 0.513834f
C530 magic_comp_0/magic_xnor_1/magic_nand_2/a_100_n230# VSS 0.028228f
C531 magic_comp_0/magic_xnor_1/magic_nand_1/Y VSS 0.570102f
C532 S1 VSS 2.942406f
C533 magic_comp_0/magic_xnor_1/magic_nand_1/a_100_n230# VSS 0.028228f
C534 magic_comp_0/magic_and_0/A VSS 1.481206f
C535 magic_comp_0/magic_xnor_1/magic_nand_0/a_100_n230# VSS 0.028228f
C536 magic_comp_0/magic_xnor_0/magic_nand_2/Y VSS 0.735888f
C537 magic_comp_0/magic_xnor_0/magic_inv_1/Y VSS 0.876873f
C538 magic_comp_0/magic_xnor_0/magic_inv_0/Y VSS 0.513834f
C539 magic_comp_0/magic_xnor_0/magic_nand_2/a_100_n230# VSS 0.028228f
C540 magic_comp_0/magic_xnor_0/magic_nand_1/Y VSS 0.570133f
C541 S0 VSS 1.962806f
C542 magic_comp_0/magic_xnor_0/magic_nand_1/a_100_n230# VSS 0.028228f
C543 magic_comp_0/magic_and_0/B VSS 1.360612f
C544 magic_comp_0/magic_xnor_0/magic_nand_0/a_100_n230# VSS 0.028228f
C545 clk VSS 13.885652f
C546 magic_dff_0/magic_nand_3/Y VSS 0.625399f
C547 magic_dff_0/magic_nand_3/a_100_n230# VSS 0.028228f
C548 magic_dff_0/magic_nand_2/Y VSS 0.673454f
C549 magic_comp_0/Y VSS 3.620044f
C550 magic_dff_0/magic_inv_0/Y VSS 0.53718f
C551 magic_dff_0/magic_nand_2/a_100_n230# VSS 0.028228f
C552 magic_dff_0/Q VSS 5.870831f
C553 magic_dff_0/magic_nand_1/a_100_n230# VSS 0.030632f
C554 magic_dff_0/notQ VSS 1.090789f
C555 magic_dff_0/magic_nand_0/a_100_n230# VSS 0.028228f
C556 magic_nand_1/A VSS 0.672088f
C557 magic_nand_1/a_100_n230# VSS 0.011246f
C558 magic_nand_0/a_100_n230# VSS 0.029249f
.ends

