** xnor.cir
.include xnor.spice
Xxnor VDD A B Y VSS xnor
.end

