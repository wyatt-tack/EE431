** xnor_magic.cir
.include magic_xnor.spice 
Xxnor A B Y VDD VSS magic_xnor
.end

