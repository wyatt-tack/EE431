magic
tech sky130A
timestamp 1731534886
<< error_p >>
rect -40 -140 -15 -138
rect -62 -160 -55 -155
rect -45 -158 -38 -140
rect -45 -160 -33 -158
rect -12 -160 0 -158
rect -45 -170 0 -168
rect -57 -185 -55 -170
rect 10 -185 12 -170
rect -45 -197 -33 -190
rect -12 -197 0 -190
<< nwell >>
rect -105 180 215 430
<< nmos >>
rect 0 -115 50 85
rect 100 -115 150 85
<< pmos >>
rect 0 200 50 400
rect 100 200 150 400
<< ndiff >>
rect -45 70 0 85
rect -45 -100 -35 70
rect -15 -100 0 70
rect -45 -115 0 -100
rect 50 30 100 85
rect 50 -110 55 30
rect 95 -110 100 30
rect 50 -115 100 -110
rect 150 70 195 85
rect 150 -100 165 70
rect 185 -100 195 70
rect 150 -115 195 -100
<< pdiff >>
rect -45 385 0 400
rect -45 215 -35 385
rect -15 215 0 385
rect -45 200 0 215
rect 50 385 100 400
rect 50 215 65 385
rect 85 215 100 385
rect 50 200 100 215
rect 150 385 195 400
rect 150 215 165 385
rect 185 215 195 385
rect 150 200 195 215
<< ndiffc >>
rect -35 -100 -15 70
rect 165 -100 185 70
<< pdiffc >>
rect -35 215 -15 385
rect 65 215 85 385
rect 165 215 185 385
<< psubdiff >>
rect -55 -170 10 -160
rect -55 -185 -45 -170
rect 0 -185 10 -170
rect -55 -190 10 -185
<< nsubdiff >>
rect -85 385 -45 400
rect -85 215 -75 385
rect -55 215 -45 385
rect -85 200 -45 215
<< psubdiffcont >>
rect -45 -185 0 -170
<< nsubdiffcont >>
rect -75 215 -55 385
<< poly >>
rect 0 400 50 415
rect 100 400 150 415
rect 0 180 50 200
rect -40 175 50 180
rect -40 155 5 175
rect 25 155 50 175
rect -40 150 50 155
rect 0 85 50 150
rect 100 125 150 200
rect 100 105 105 125
rect 125 105 150 125
rect 100 85 150 105
rect 0 -130 50 -115
rect 100 -130 150 -115
<< polycont >>
rect 5 155 25 175
rect 105 105 125 125
<< ndiffres >>
rect 55 -110 95 30
<< locali >>
rect -85 425 -65 430
rect -85 390 -65 405
rect 155 425 175 430
rect 155 390 175 405
rect -85 385 -5 390
rect -85 215 -75 385
rect -55 215 -35 385
rect -15 215 -5 385
rect -85 210 -5 215
rect 55 385 95 390
rect 55 215 65 385
rect 85 215 95 385
rect 55 180 95 215
rect 155 385 195 390
rect 155 215 165 385
rect 185 215 195 385
rect 155 210 195 215
rect -105 175 35 180
rect -105 155 5 175
rect 25 155 35 175
rect -105 150 35 155
rect 55 150 215 180
rect -105 125 135 130
rect -105 105 105 125
rect 125 105 135 125
rect -105 100 135 105
rect -45 70 -5 75
rect -45 -100 -35 70
rect -15 -100 -5 70
rect -85 -135 -65 -130
rect -45 -140 -5 -100
rect 155 70 195 150
rect 155 -100 165 70
rect 185 -100 195 70
rect 155 -115 195 -100
rect -45 -155 -40 -140
rect -15 -155 -5 -140
rect -85 -160 -55 -155
rect -45 -160 -5 -155
rect -85 -170 10 -160
rect -85 -185 -45 -170
rect 0 -185 10 -170
rect -85 -190 10 -185
<< viali >>
rect -85 405 -65 425
rect 155 405 175 425
rect -85 -155 -65 -135
rect -40 -155 -15 -140
<< metal1 >>
rect -105 425 215 430
rect -105 405 -85 425
rect -65 405 155 425
rect 175 405 215 425
rect -105 400 215 405
rect -105 -135 220 -130
rect -105 -155 -85 -135
rect -65 -140 220 -135
rect -65 -155 -40 -140
rect -15 -155 220 -140
rect -105 -160 220 -155
<< labels >>
rlabel locali -105 150 -85 180 7 A
port 1 w
rlabel locali -105 100 -85 130 7 B
port 2 w
rlabel locali 195 150 215 180 3 Y
port 3 e
rlabel metal1 -105 400 -85 430 7 VDD
port 4 w
rlabel metal1 -105 -160 -85 -130 7 VSS
port 5 w
<< end >>
