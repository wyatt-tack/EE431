magic
tech sky130A
timestamp 1733267924
<< nwell >>
rect 5950 665 6155 915
<< poly >>
rect -70 2555 255 2560
rect -70 2535 -60 2555
rect -40 2535 255 2555
rect -70 2530 255 2535
rect -70 -1585 -40 2530
rect 5685 2475 8080 2510
rect 5685 1945 5715 2475
rect 8030 2435 8080 2475
rect 5685 1925 5690 1945
rect 5710 1925 5715 1945
rect 5685 1915 5715 1925
rect 5790 225 5840 370
rect 5610 195 5840 225
rect 5890 225 5940 370
rect 5890 195 8005 225
rect 5340 -20 5370 -10
rect 15 -25 1995 -20
rect 15 -45 1965 -25
rect 1985 -45 1995 -25
rect 15 -50 1995 -45
rect 5340 -40 5345 -20
rect 5365 -40 5370 -20
rect 15 -510 45 -50
rect 5 -515 45 -510
rect 5 -535 15 -515
rect 35 -535 45 -515
rect 5 -540 45 -535
rect 70 -80 1995 -75
rect 70 -100 1965 -80
rect 1985 -100 1995 -80
rect 70 -105 1995 -100
rect 70 -560 100 -105
rect 60 -565 100 -560
rect 60 -585 70 -565
rect 90 -585 100 -565
rect 60 -590 100 -585
rect 125 -135 1995 -130
rect 125 -155 1965 -135
rect 1985 -155 1995 -135
rect 125 -160 1995 -155
rect 125 -610 155 -160
rect 115 -615 155 -610
rect 115 -635 125 -615
rect 145 -635 155 -615
rect 115 -640 155 -635
rect 180 -190 1995 -185
rect 180 -210 1965 -190
rect 1985 -210 1995 -190
rect 180 -215 1995 -210
rect 180 -660 210 -215
rect 170 -665 210 -660
rect 170 -685 180 -665
rect 200 -685 210 -665
rect 170 -690 210 -685
rect 4235 -310 4265 -300
rect 4235 -330 4240 -310
rect 4260 -330 4265 -310
rect 4235 -1260 4265 -330
rect 5340 -335 5370 -40
rect 5610 -335 5650 195
rect 7955 90 8005 195
rect 5340 -340 5650 -335
rect 5340 -360 5620 -340
rect 5640 -360 5650 -340
rect 5340 -365 5650 -360
rect 7000 50 7030 60
rect 7000 30 7005 50
rect 7025 30 7030 50
rect 7000 -1175 7030 30
rect 5475 -1180 7030 -1175
rect 5475 -1200 5485 -1180
rect 5505 -1200 7030 -1180
rect 5475 -1205 7030 -1200
rect 4235 -1265 4275 -1260
rect 4235 -1285 4245 -1265
rect 4265 -1285 4275 -1265
rect 4235 -1290 4275 -1285
rect 4235 -1585 4265 -1290
rect -70 -1615 4265 -1585
<< polycont >>
rect -60 2535 -40 2555
rect 5690 1925 5710 1945
rect 1965 -45 1985 -25
rect 5345 -40 5365 -20
rect 15 -535 35 -515
rect 1965 -100 1985 -80
rect 70 -585 90 -565
rect 1965 -155 1985 -135
rect 125 -635 145 -615
rect 1965 -210 1985 -190
rect 180 -685 200 -665
rect 4240 -330 4260 -310
rect 5620 -360 5640 -340
rect 7005 30 7025 50
rect 5485 -1200 5505 -1180
rect 4245 -1285 4265 -1265
<< locali >>
rect 5420 2590 5570 2620
rect -125 2555 255 2560
rect -125 2535 -60 2555
rect -40 2535 255 2555
rect -125 2530 255 2535
rect 5415 2530 5520 2560
rect 5405 1375 5470 1405
rect 5340 -20 5370 1095
rect 1955 -25 5345 -20
rect 1955 -45 1965 -25
rect 1985 -40 5345 -25
rect 5365 -40 5370 -20
rect 1985 -45 5370 -40
rect 1955 -50 5370 -45
rect 5440 -75 5470 1375
rect 1955 -80 5470 -75
rect 1955 -100 1965 -80
rect 1985 -100 5470 -80
rect 1955 -105 5470 -100
rect 5490 -130 5520 2530
rect 1955 -135 5520 -130
rect 1955 -155 1965 -135
rect 1985 -155 5520 -135
rect 1955 -160 5520 -155
rect 5540 -185 5570 2590
rect 5610 2170 5690 2200
rect 8235 2170 8280 2200
rect 5610 1035 5640 2170
rect 5685 1945 5715 1955
rect 5685 1925 5690 1945
rect 5710 1925 5715 1945
rect 5685 1915 5715 1925
rect 5610 995 6290 1035
rect 6250 825 6290 995
rect 5955 635 6150 665
rect 6255 265 6285 615
rect 6255 235 7030 265
rect 7000 50 7030 235
rect 7000 30 7005 50
rect 7025 30 7030 50
rect 7000 20 7030 30
rect 1955 -190 5570 -185
rect 1955 -210 1965 -190
rect 1985 -210 5570 -190
rect 1955 -215 5570 -210
rect 5610 -270 5640 -80
rect 4235 -300 5640 -270
rect 4235 -310 4265 -300
rect 4235 -330 4240 -310
rect 4260 -330 4265 -310
rect 4235 -340 4265 -330
rect 5 -515 180 -510
rect 5 -535 15 -515
rect 35 -535 180 -515
rect 5 -540 180 -535
rect 60 -565 180 -560
rect 60 -585 70 -565
rect 90 -585 180 -565
rect 60 -590 180 -585
rect 115 -615 180 -610
rect 115 -635 125 -615
rect 145 -635 180 -615
rect 115 -640 180 -635
rect 170 -690 180 -660
rect -125 -760 200 -730
rect -125 -815 200 -785
rect -125 -870 200 -840
rect -125 -925 200 -895
rect 5475 -1180 5515 -1175
rect 5475 -1200 5485 -1180
rect 5505 -1200 5515 -1180
rect 5475 -1205 5515 -1200
rect 4185 -1240 4455 -1210
rect 5205 -1240 5515 -1205
rect 4185 -1910 4215 -1240
rect 4235 -1265 4350 -1260
rect 4235 -1285 4245 -1265
rect 4265 -1285 4350 -1265
rect 4235 -1290 4350 -1285
<< metal1 >>
rect -125 2785 8280 2840
rect -125 2780 95 2785
rect 5330 2780 8280 2785
rect 5260 2150 5280 2780
rect 5330 1415 5440 2780
rect 6245 2420 6295 2780
rect 5370 1365 5440 1415
rect 5330 1315 5440 1365
rect 5370 980 5440 1315
rect 8210 1150 8250 1220
rect 5370 915 5580 980
rect 5370 910 5690 915
rect 5510 885 5690 910
rect 6000 885 6100 915
rect 5510 170 5580 885
rect 6480 355 6520 1120
rect 6010 325 6110 355
rect 6400 325 6520 355
rect 5510 140 5620 170
rect 0 -2190 40 70
rect 5510 -240 5580 140
rect 4180 -270 5580 -240
rect 4350 -990 4390 -270
rect 5610 -2190 5660 -1060
rect 8200 -2190 8250 1150
rect -125 -2245 8280 -2190
use magic_comp  magic_comp_0
timestamp 1733183236
transform 1 0 335 0 1 -1570
box -155 -650 3850 1330
use magic_counter  magic_counter_0
timestamp 1732472291
transform 1 0 80 0 1 1480
box -80 -1480 5340 1330
use magic_dff  magic_dff_0
timestamp 1732136480
transform 1 0 5045 0 1 -1550
box -695 -670 390 590
use magic_etdff  magic_etdff_0
timestamp 1732138536
transform 1 0 6620 0 1 -480
box -1010 -680 1540 650
use magic_etdff  magic_etdff_1
timestamp 1732138536
transform 1 0 6695 0 1 1800
box -1010 -680 1540 650
use magic_nand  magic_nand_0
timestamp 1731535207
transform 1 0 5790 0 1 485
box -105 -160 220 430
use magic_nand  magic_nand_1
timestamp 1731535207
transform 1 0 6195 0 1 485
box -105 -160 220 430
<< labels >>
rlabel locali -125 -925 -105 -895 7 S0
port 2 w
rlabel locali -125 -870 -105 -840 7 S1
port 3 w
rlabel locali -125 -815 -105 -785 7 S2
port 4 w
rlabel locali -125 -760 -105 -730 7 S3
port 5 w
rlabel metal1 -125 2780 -105 2840 7 VDD
port 7 w
rlabel metal1 -125 -2245 -105 -2190 7 VSS
port 8 w
rlabel locali -125 2530 -105 2560 7 clk
port 1 w
rlabel locali 8260 2170 8280 2200 3 PWM
port 6 e
<< end >>
