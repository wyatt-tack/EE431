magic
tech sky130A
timestamp 1732472291
<< poly >>
rect 5280 1130 5310 1140
rect 5280 1110 5285 1130
rect 5305 1110 5310 1130
rect 2680 1050 2805 1080
rect 2680 -10 2710 1050
rect 5280 -10 5310 1110
rect 2680 -40 5310 -10
rect 2680 -80 5330 -75
rect 2680 -100 5300 -80
rect 5320 -100 5330 -80
rect 2680 -105 5330 -100
rect 2680 -365 2710 -105
rect 2680 -395 2845 -365
<< polycont >>
rect 5285 1110 5305 1130
rect 5300 -100 5320 -80
<< locali >>
rect 5280 1130 5340 1140
rect 5280 1110 5285 1130
rect 5305 1110 5340 1130
rect 5280 1100 5310 1110
rect -80 1050 0 1080
rect 2540 1050 2670 1080
rect 5215 1050 5340 1080
rect 0 0 30 825
rect 2510 0 2550 410
rect 0 -30 2550 0
rect 2680 0 2710 795
rect 5180 0 5220 410
rect 2680 -30 5220 0
rect 5240 -50 5270 1050
rect 0 -80 5270 -50
rect 5290 -80 5340 -75
rect 0 -395 30 -80
rect 5290 -100 5300 -80
rect 5320 -100 5340 -80
rect 5290 -105 5340 -100
rect 2550 -395 2680 -365
rect 5220 -395 5340 -365
rect 0 -1450 30 -620
rect 2520 -1450 2550 -1035
rect 0 -1480 2550 -1450
rect 2670 -1450 2700 -620
rect 5190 -1450 5220 -1035
rect 2670 -1480 5220 -1450
<< metal1 >>
rect -80 1300 15 1330
rect 2550 1300 2680 1330
rect 5220 1300 5340 1330
rect -80 1290 0 1300
rect 5180 630 5290 670
rect -60 0 45 40
rect 2550 0 2670 30
rect -60 -560 -20 0
rect 5250 -115 5290 630
rect 2550 -145 2680 -115
rect 5155 -165 5290 -115
rect -60 -600 45 -560
rect 20 -1410 85 -1405
rect -80 -1420 85 -1410
rect 2530 -1415 2690 -1345
rect 2545 -1420 2675 -1415
rect 5200 -1420 5220 -1345
rect -80 -1480 5340 -1420
use magic_etdff  magic_etdff_0
timestamp 1732138536
transform 1 0 1010 0 1 680
box -1010 -680 1540 650
use magic_etdff  magic_etdff_1
timestamp 1732138536
transform 1 0 3680 0 1 680
box -1010 -680 1540 650
use magic_etdff  magic_etdff_2
timestamp 1732138536
transform 1 0 1010 0 1 -765
box -1010 -680 1540 650
use magic_etdff  magic_etdff_3
timestamp 1732138536
transform 1 0 3680 0 1 -765
box -1010 -680 1540 650
<< labels >>
rlabel locali -80 1050 -60 1080 7 clk
port 1 w
rlabel locali 5320 -105 5340 -75 3 S2
port 4 e
rlabel locali 5320 -395 5340 -365 3 S3
port 5 e
rlabel metal1 -80 1290 -60 1330 7 VDD
port 6 w
rlabel metal1 -80 -1480 -60 -1410 7 VSS
port 7 w
rlabel locali 5320 1110 5340 1140 3 S0
port 2 e
rlabel locali 5320 1050 5340 1080 3 S1
port 3 e
<< end >>
