** inv_magic.cir
.include magic_nand.spice
Xnand A B Y VDD VSS magic_nand
.end

