magic
tech sky130A
timestamp 1732493268
<< poly >>
rect -5 -30 1970 0
rect -5 -85 1370 -55
rect -5 -140 780 -110
rect -5 -195 140 -165
rect 110 -200 140 -195
rect 750 -200 780 -140
rect 1340 -200 1370 -85
rect 1940 -200 1970 -30
<< locali >>
rect 5420 2590 5570 2620
rect 5415 2530 5520 2560
rect 5405 1375 5470 1405
rect 5340 -20 5370 1095
rect 120 -50 5370 -20
rect 120 -200 150 -50
rect 5440 -70 5470 1375
rect 730 -200 750 -70
rect 5395 -100 5470 -70
rect 5490 -120 5520 2530
rect 1330 -150 5520 -120
rect 1330 -200 1350 -150
rect 5540 -170 5570 2590
rect 1930 -200 1950 -170
rect 5460 -200 5570 -170
<< rlocali >>
rect 750 -100 5395 -70
rect 1950 -200 5460 -170
<< metal1 >>
rect 5370 1365 5440 1415
rect 5330 1315 5440 1365
rect 5370 980 5440 1315
rect 5370 910 5580 980
rect 5510 -200 5580 910
use magic_counter  magic_counter_0
timestamp 1732472291
transform 1 0 80 0 1 1480
box -80 -1480 5340 1330
<< end >>
